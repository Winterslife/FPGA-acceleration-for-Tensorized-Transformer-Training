
    wire dl_reset;
    wire dl_clock;
    assign dl_reset = ap_rst_n;
    assign dl_clock = ap_clk;
    wire [33:0] proc_0_data_FIFO_blk;
    wire [33:0] proc_0_data_PIPO_blk;
    wire [33:0] proc_0_start_FIFO_blk;
    wire [33:0] proc_0_TLF_FIFO_blk;
    wire [33:0] proc_0_input_sync_blk;
    wire [33:0] proc_0_output_sync_blk;
    wire [33:0] proc_dep_vld_vec_0;
    reg [33:0] proc_dep_vld_vec_0_reg;
    wire [33:0] in_chan_dep_vld_vec_0;
    wire [1359:0] in_chan_dep_data_vec_0;
    wire [33:0] token_in_vec_0;
    wire [33:0] out_chan_dep_vld_vec_0;
    wire [39:0] out_chan_dep_data_0;
    wire [33:0] token_out_vec_0;
    wire dl_detect_out_0;
    wire dep_chan_vld_1_0;
    wire [39:0] dep_chan_data_1_0;
    wire token_1_0;
    wire dep_chan_vld_3_0;
    wire [39:0] dep_chan_data_3_0;
    wire token_3_0;
    wire dep_chan_vld_6_0;
    wire [39:0] dep_chan_data_6_0;
    wire token_6_0;
    wire dep_chan_vld_7_0;
    wire [39:0] dep_chan_data_7_0;
    wire token_7_0;
    wire dep_chan_vld_8_0;
    wire [39:0] dep_chan_data_8_0;
    wire token_8_0;
    wire dep_chan_vld_9_0;
    wire [39:0] dep_chan_data_9_0;
    wire token_9_0;
    wire dep_chan_vld_10_0;
    wire [39:0] dep_chan_data_10_0;
    wire token_10_0;
    wire dep_chan_vld_11_0;
    wire [39:0] dep_chan_data_11_0;
    wire token_11_0;
    wire dep_chan_vld_12_0;
    wire [39:0] dep_chan_data_12_0;
    wire token_12_0;
    wire dep_chan_vld_13_0;
    wire [39:0] dep_chan_data_13_0;
    wire token_13_0;
    wire dep_chan_vld_14_0;
    wire [39:0] dep_chan_data_14_0;
    wire token_14_0;
    wire dep_chan_vld_15_0;
    wire [39:0] dep_chan_data_15_0;
    wire token_15_0;
    wire dep_chan_vld_16_0;
    wire [39:0] dep_chan_data_16_0;
    wire token_16_0;
    wire dep_chan_vld_17_0;
    wire [39:0] dep_chan_data_17_0;
    wire token_17_0;
    wire dep_chan_vld_18_0;
    wire [39:0] dep_chan_data_18_0;
    wire token_18_0;
    wire dep_chan_vld_19_0;
    wire [39:0] dep_chan_data_19_0;
    wire token_19_0;
    wire dep_chan_vld_20_0;
    wire [39:0] dep_chan_data_20_0;
    wire token_20_0;
    wire dep_chan_vld_21_0;
    wire [39:0] dep_chan_data_21_0;
    wire token_21_0;
    wire dep_chan_vld_22_0;
    wire [39:0] dep_chan_data_22_0;
    wire token_22_0;
    wire dep_chan_vld_23_0;
    wire [39:0] dep_chan_data_23_0;
    wire token_23_0;
    wire dep_chan_vld_24_0;
    wire [39:0] dep_chan_data_24_0;
    wire token_24_0;
    wire dep_chan_vld_25_0;
    wire [39:0] dep_chan_data_25_0;
    wire token_25_0;
    wire dep_chan_vld_26_0;
    wire [39:0] dep_chan_data_26_0;
    wire token_26_0;
    wire dep_chan_vld_27_0;
    wire [39:0] dep_chan_data_27_0;
    wire token_27_0;
    wire dep_chan_vld_28_0;
    wire [39:0] dep_chan_data_28_0;
    wire token_28_0;
    wire dep_chan_vld_29_0;
    wire [39:0] dep_chan_data_29_0;
    wire token_29_0;
    wire dep_chan_vld_30_0;
    wire [39:0] dep_chan_data_30_0;
    wire token_30_0;
    wire dep_chan_vld_31_0;
    wire [39:0] dep_chan_data_31_0;
    wire token_31_0;
    wire dep_chan_vld_32_0;
    wire [39:0] dep_chan_data_32_0;
    wire token_32_0;
    wire dep_chan_vld_33_0;
    wire [39:0] dep_chan_data_33_0;
    wire token_33_0;
    wire dep_chan_vld_34_0;
    wire [39:0] dep_chan_data_34_0;
    wire token_34_0;
    wire dep_chan_vld_35_0;
    wire [39:0] dep_chan_data_35_0;
    wire token_35_0;
    wire dep_chan_vld_36_0;
    wire [39:0] dep_chan_data_36_0;
    wire token_36_0;
    wire dep_chan_vld_39_0;
    wire [39:0] dep_chan_data_39_0;
    wire token_39_0;
    wire [33:0] proc_1_data_FIFO_blk;
    wire [33:0] proc_1_data_PIPO_blk;
    wire [33:0] proc_1_start_FIFO_blk;
    wire [33:0] proc_1_TLF_FIFO_blk;
    wire [33:0] proc_1_input_sync_blk;
    wire [33:0] proc_1_output_sync_blk;
    wire [33:0] proc_dep_vld_vec_1;
    reg [33:0] proc_dep_vld_vec_1_reg;
    wire [33:0] in_chan_dep_vld_vec_1;
    wire [1359:0] in_chan_dep_data_vec_1;
    wire [33:0] token_in_vec_1;
    wire [33:0] out_chan_dep_vld_vec_1;
    wire [39:0] out_chan_dep_data_1;
    wire [33:0] token_out_vec_1;
    wire dl_detect_out_1;
    wire dep_chan_vld_0_1;
    wire [39:0] dep_chan_data_0_1;
    wire token_0_1;
    wire dep_chan_vld_2_1;
    wire [39:0] dep_chan_data_2_1;
    wire token_2_1;
    wire dep_chan_vld_3_1;
    wire [39:0] dep_chan_data_3_1;
    wire token_3_1;
    wire dep_chan_vld_6_1;
    wire [39:0] dep_chan_data_6_1;
    wire token_6_1;
    wire dep_chan_vld_7_1;
    wire [39:0] dep_chan_data_7_1;
    wire token_7_1;
    wire dep_chan_vld_8_1;
    wire [39:0] dep_chan_data_8_1;
    wire token_8_1;
    wire dep_chan_vld_9_1;
    wire [39:0] dep_chan_data_9_1;
    wire token_9_1;
    wire dep_chan_vld_10_1;
    wire [39:0] dep_chan_data_10_1;
    wire token_10_1;
    wire dep_chan_vld_11_1;
    wire [39:0] dep_chan_data_11_1;
    wire token_11_1;
    wire dep_chan_vld_12_1;
    wire [39:0] dep_chan_data_12_1;
    wire token_12_1;
    wire dep_chan_vld_13_1;
    wire [39:0] dep_chan_data_13_1;
    wire token_13_1;
    wire dep_chan_vld_14_1;
    wire [39:0] dep_chan_data_14_1;
    wire token_14_1;
    wire dep_chan_vld_15_1;
    wire [39:0] dep_chan_data_15_1;
    wire token_15_1;
    wire dep_chan_vld_16_1;
    wire [39:0] dep_chan_data_16_1;
    wire token_16_1;
    wire dep_chan_vld_17_1;
    wire [39:0] dep_chan_data_17_1;
    wire token_17_1;
    wire dep_chan_vld_18_1;
    wire [39:0] dep_chan_data_18_1;
    wire token_18_1;
    wire dep_chan_vld_19_1;
    wire [39:0] dep_chan_data_19_1;
    wire token_19_1;
    wire dep_chan_vld_20_1;
    wire [39:0] dep_chan_data_20_1;
    wire token_20_1;
    wire dep_chan_vld_21_1;
    wire [39:0] dep_chan_data_21_1;
    wire token_21_1;
    wire dep_chan_vld_22_1;
    wire [39:0] dep_chan_data_22_1;
    wire token_22_1;
    wire dep_chan_vld_23_1;
    wire [39:0] dep_chan_data_23_1;
    wire token_23_1;
    wire dep_chan_vld_24_1;
    wire [39:0] dep_chan_data_24_1;
    wire token_24_1;
    wire dep_chan_vld_25_1;
    wire [39:0] dep_chan_data_25_1;
    wire token_25_1;
    wire dep_chan_vld_26_1;
    wire [39:0] dep_chan_data_26_1;
    wire token_26_1;
    wire dep_chan_vld_27_1;
    wire [39:0] dep_chan_data_27_1;
    wire token_27_1;
    wire dep_chan_vld_28_1;
    wire [39:0] dep_chan_data_28_1;
    wire token_28_1;
    wire dep_chan_vld_29_1;
    wire [39:0] dep_chan_data_29_1;
    wire token_29_1;
    wire dep_chan_vld_30_1;
    wire [39:0] dep_chan_data_30_1;
    wire token_30_1;
    wire dep_chan_vld_31_1;
    wire [39:0] dep_chan_data_31_1;
    wire token_31_1;
    wire dep_chan_vld_32_1;
    wire [39:0] dep_chan_data_32_1;
    wire token_32_1;
    wire dep_chan_vld_33_1;
    wire [39:0] dep_chan_data_33_1;
    wire token_33_1;
    wire dep_chan_vld_34_1;
    wire [39:0] dep_chan_data_34_1;
    wire token_34_1;
    wire dep_chan_vld_35_1;
    wire [39:0] dep_chan_data_35_1;
    wire token_35_1;
    wire dep_chan_vld_36_1;
    wire [39:0] dep_chan_data_36_1;
    wire token_36_1;
    wire [1:0] proc_2_data_FIFO_blk;
    wire [1:0] proc_2_data_PIPO_blk;
    wire [1:0] proc_2_start_FIFO_blk;
    wire [1:0] proc_2_TLF_FIFO_blk;
    wire [1:0] proc_2_input_sync_blk;
    wire [1:0] proc_2_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_2;
    reg [1:0] proc_dep_vld_vec_2_reg;
    wire [1:0] in_chan_dep_vld_vec_2;
    wire [79:0] in_chan_dep_data_vec_2;
    wire [1:0] token_in_vec_2;
    wire [1:0] out_chan_dep_vld_vec_2;
    wire [39:0] out_chan_dep_data_2;
    wire [1:0] token_out_vec_2;
    wire dl_detect_out_2;
    wire dep_chan_vld_1_2;
    wire [39:0] dep_chan_data_1_2;
    wire token_1_2;
    wire dep_chan_vld_6_2;
    wire [39:0] dep_chan_data_6_2;
    wire token_6_2;
    wire [33:0] proc_3_data_FIFO_blk;
    wire [33:0] proc_3_data_PIPO_blk;
    wire [33:0] proc_3_start_FIFO_blk;
    wire [33:0] proc_3_TLF_FIFO_blk;
    wire [33:0] proc_3_input_sync_blk;
    wire [33:0] proc_3_output_sync_blk;
    wire [33:0] proc_dep_vld_vec_3;
    reg [33:0] proc_dep_vld_vec_3_reg;
    wire [33:0] in_chan_dep_vld_vec_3;
    wire [1359:0] in_chan_dep_data_vec_3;
    wire [33:0] token_in_vec_3;
    wire [33:0] out_chan_dep_vld_vec_3;
    wire [39:0] out_chan_dep_data_3;
    wire [33:0] token_out_vec_3;
    wire dl_detect_out_3;
    wire dep_chan_vld_0_3;
    wire [39:0] dep_chan_data_0_3;
    wire token_0_3;
    wire dep_chan_vld_1_3;
    wire [39:0] dep_chan_data_1_3;
    wire token_1_3;
    wire dep_chan_vld_4_3;
    wire [39:0] dep_chan_data_4_3;
    wire token_4_3;
    wire dep_chan_vld_6_3;
    wire [39:0] dep_chan_data_6_3;
    wire token_6_3;
    wire dep_chan_vld_7_3;
    wire [39:0] dep_chan_data_7_3;
    wire token_7_3;
    wire dep_chan_vld_8_3;
    wire [39:0] dep_chan_data_8_3;
    wire token_8_3;
    wire dep_chan_vld_9_3;
    wire [39:0] dep_chan_data_9_3;
    wire token_9_3;
    wire dep_chan_vld_10_3;
    wire [39:0] dep_chan_data_10_3;
    wire token_10_3;
    wire dep_chan_vld_11_3;
    wire [39:0] dep_chan_data_11_3;
    wire token_11_3;
    wire dep_chan_vld_12_3;
    wire [39:0] dep_chan_data_12_3;
    wire token_12_3;
    wire dep_chan_vld_13_3;
    wire [39:0] dep_chan_data_13_3;
    wire token_13_3;
    wire dep_chan_vld_14_3;
    wire [39:0] dep_chan_data_14_3;
    wire token_14_3;
    wire dep_chan_vld_15_3;
    wire [39:0] dep_chan_data_15_3;
    wire token_15_3;
    wire dep_chan_vld_16_3;
    wire [39:0] dep_chan_data_16_3;
    wire token_16_3;
    wire dep_chan_vld_17_3;
    wire [39:0] dep_chan_data_17_3;
    wire token_17_3;
    wire dep_chan_vld_18_3;
    wire [39:0] dep_chan_data_18_3;
    wire token_18_3;
    wire dep_chan_vld_19_3;
    wire [39:0] dep_chan_data_19_3;
    wire token_19_3;
    wire dep_chan_vld_20_3;
    wire [39:0] dep_chan_data_20_3;
    wire token_20_3;
    wire dep_chan_vld_21_3;
    wire [39:0] dep_chan_data_21_3;
    wire token_21_3;
    wire dep_chan_vld_22_3;
    wire [39:0] dep_chan_data_22_3;
    wire token_22_3;
    wire dep_chan_vld_23_3;
    wire [39:0] dep_chan_data_23_3;
    wire token_23_3;
    wire dep_chan_vld_24_3;
    wire [39:0] dep_chan_data_24_3;
    wire token_24_3;
    wire dep_chan_vld_25_3;
    wire [39:0] dep_chan_data_25_3;
    wire token_25_3;
    wire dep_chan_vld_26_3;
    wire [39:0] dep_chan_data_26_3;
    wire token_26_3;
    wire dep_chan_vld_27_3;
    wire [39:0] dep_chan_data_27_3;
    wire token_27_3;
    wire dep_chan_vld_28_3;
    wire [39:0] dep_chan_data_28_3;
    wire token_28_3;
    wire dep_chan_vld_29_3;
    wire [39:0] dep_chan_data_29_3;
    wire token_29_3;
    wire dep_chan_vld_30_3;
    wire [39:0] dep_chan_data_30_3;
    wire token_30_3;
    wire dep_chan_vld_31_3;
    wire [39:0] dep_chan_data_31_3;
    wire token_31_3;
    wire dep_chan_vld_32_3;
    wire [39:0] dep_chan_data_32_3;
    wire token_32_3;
    wire dep_chan_vld_33_3;
    wire [39:0] dep_chan_data_33_3;
    wire token_33_3;
    wire dep_chan_vld_34_3;
    wire [39:0] dep_chan_data_34_3;
    wire token_34_3;
    wire dep_chan_vld_35_3;
    wire [39:0] dep_chan_data_35_3;
    wire token_35_3;
    wire dep_chan_vld_36_3;
    wire [39:0] dep_chan_data_36_3;
    wire token_36_3;
    wire [1:0] proc_4_data_FIFO_blk;
    wire [1:0] proc_4_data_PIPO_blk;
    wire [1:0] proc_4_start_FIFO_blk;
    wire [1:0] proc_4_TLF_FIFO_blk;
    wire [1:0] proc_4_input_sync_blk;
    wire [1:0] proc_4_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_4;
    reg [1:0] proc_dep_vld_vec_4_reg;
    wire [1:0] in_chan_dep_vld_vec_4;
    wire [79:0] in_chan_dep_data_vec_4;
    wire [1:0] token_in_vec_4;
    wire [1:0] out_chan_dep_vld_vec_4;
    wire [39:0] out_chan_dep_data_4;
    wire [1:0] token_out_vec_4;
    wire dl_detect_out_4;
    wire dep_chan_vld_3_4;
    wire [39:0] dep_chan_data_3_4;
    wire token_3_4;
    wire dep_chan_vld_5_4;
    wire [39:0] dep_chan_data_5_4;
    wire token_5_4;
    wire [1:0] proc_5_data_FIFO_blk;
    wire [1:0] proc_5_data_PIPO_blk;
    wire [1:0] proc_5_start_FIFO_blk;
    wire [1:0] proc_5_TLF_FIFO_blk;
    wire [1:0] proc_5_input_sync_blk;
    wire [1:0] proc_5_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_5;
    reg [1:0] proc_dep_vld_vec_5_reg;
    wire [1:0] in_chan_dep_vld_vec_5;
    wire [79:0] in_chan_dep_data_vec_5;
    wire [1:0] token_in_vec_5;
    wire [1:0] out_chan_dep_vld_vec_5;
    wire [39:0] out_chan_dep_data_5;
    wire [1:0] token_out_vec_5;
    wire dl_detect_out_5;
    wire dep_chan_vld_4_5;
    wire [39:0] dep_chan_data_4_5;
    wire token_4_5;
    wire dep_chan_vld_6_5;
    wire [39:0] dep_chan_data_6_5;
    wire token_6_5;
    wire [35:0] proc_6_data_FIFO_blk;
    wire [35:0] proc_6_data_PIPO_blk;
    wire [35:0] proc_6_start_FIFO_blk;
    wire [35:0] proc_6_TLF_FIFO_blk;
    wire [35:0] proc_6_input_sync_blk;
    wire [35:0] proc_6_output_sync_blk;
    wire [35:0] proc_dep_vld_vec_6;
    reg [35:0] proc_dep_vld_vec_6_reg;
    wire [35:0] in_chan_dep_vld_vec_6;
    wire [1439:0] in_chan_dep_data_vec_6;
    wire [35:0] token_in_vec_6;
    wire [35:0] out_chan_dep_vld_vec_6;
    wire [39:0] out_chan_dep_data_6;
    wire [35:0] token_out_vec_6;
    wire dl_detect_out_6;
    wire dep_chan_vld_0_6;
    wire [39:0] dep_chan_data_0_6;
    wire token_0_6;
    wire dep_chan_vld_1_6;
    wire [39:0] dep_chan_data_1_6;
    wire token_1_6;
    wire dep_chan_vld_2_6;
    wire [39:0] dep_chan_data_2_6;
    wire token_2_6;
    wire dep_chan_vld_3_6;
    wire [39:0] dep_chan_data_3_6;
    wire token_3_6;
    wire dep_chan_vld_5_6;
    wire [39:0] dep_chan_data_5_6;
    wire token_5_6;
    wire dep_chan_vld_7_6;
    wire [39:0] dep_chan_data_7_6;
    wire token_7_6;
    wire dep_chan_vld_8_6;
    wire [39:0] dep_chan_data_8_6;
    wire token_8_6;
    wire dep_chan_vld_9_6;
    wire [39:0] dep_chan_data_9_6;
    wire token_9_6;
    wire dep_chan_vld_10_6;
    wire [39:0] dep_chan_data_10_6;
    wire token_10_6;
    wire dep_chan_vld_11_6;
    wire [39:0] dep_chan_data_11_6;
    wire token_11_6;
    wire dep_chan_vld_12_6;
    wire [39:0] dep_chan_data_12_6;
    wire token_12_6;
    wire dep_chan_vld_13_6;
    wire [39:0] dep_chan_data_13_6;
    wire token_13_6;
    wire dep_chan_vld_14_6;
    wire [39:0] dep_chan_data_14_6;
    wire token_14_6;
    wire dep_chan_vld_15_6;
    wire [39:0] dep_chan_data_15_6;
    wire token_15_6;
    wire dep_chan_vld_16_6;
    wire [39:0] dep_chan_data_16_6;
    wire token_16_6;
    wire dep_chan_vld_17_6;
    wire [39:0] dep_chan_data_17_6;
    wire token_17_6;
    wire dep_chan_vld_18_6;
    wire [39:0] dep_chan_data_18_6;
    wire token_18_6;
    wire dep_chan_vld_19_6;
    wire [39:0] dep_chan_data_19_6;
    wire token_19_6;
    wire dep_chan_vld_20_6;
    wire [39:0] dep_chan_data_20_6;
    wire token_20_6;
    wire dep_chan_vld_21_6;
    wire [39:0] dep_chan_data_21_6;
    wire token_21_6;
    wire dep_chan_vld_22_6;
    wire [39:0] dep_chan_data_22_6;
    wire token_22_6;
    wire dep_chan_vld_23_6;
    wire [39:0] dep_chan_data_23_6;
    wire token_23_6;
    wire dep_chan_vld_24_6;
    wire [39:0] dep_chan_data_24_6;
    wire token_24_6;
    wire dep_chan_vld_25_6;
    wire [39:0] dep_chan_data_25_6;
    wire token_25_6;
    wire dep_chan_vld_26_6;
    wire [39:0] dep_chan_data_26_6;
    wire token_26_6;
    wire dep_chan_vld_27_6;
    wire [39:0] dep_chan_data_27_6;
    wire token_27_6;
    wire dep_chan_vld_28_6;
    wire [39:0] dep_chan_data_28_6;
    wire token_28_6;
    wire dep_chan_vld_29_6;
    wire [39:0] dep_chan_data_29_6;
    wire token_29_6;
    wire dep_chan_vld_30_6;
    wire [39:0] dep_chan_data_30_6;
    wire token_30_6;
    wire dep_chan_vld_31_6;
    wire [39:0] dep_chan_data_31_6;
    wire token_31_6;
    wire dep_chan_vld_32_6;
    wire [39:0] dep_chan_data_32_6;
    wire token_32_6;
    wire dep_chan_vld_33_6;
    wire [39:0] dep_chan_data_33_6;
    wire token_33_6;
    wire dep_chan_vld_34_6;
    wire [39:0] dep_chan_data_34_6;
    wire token_34_6;
    wire dep_chan_vld_35_6;
    wire [39:0] dep_chan_data_35_6;
    wire token_35_6;
    wire dep_chan_vld_36_6;
    wire [39:0] dep_chan_data_36_6;
    wire token_36_6;
    wire dep_chan_vld_38_6;
    wire [39:0] dep_chan_data_38_6;
    wire token_38_6;
    wire [32:0] proc_7_data_FIFO_blk;
    wire [32:0] proc_7_data_PIPO_blk;
    wire [32:0] proc_7_start_FIFO_blk;
    wire [32:0] proc_7_TLF_FIFO_blk;
    wire [32:0] proc_7_input_sync_blk;
    wire [32:0] proc_7_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_7;
    reg [32:0] proc_dep_vld_vec_7_reg;
    wire [32:0] in_chan_dep_vld_vec_7;
    wire [1319:0] in_chan_dep_data_vec_7;
    wire [32:0] token_in_vec_7;
    wire [32:0] out_chan_dep_vld_vec_7;
    wire [39:0] out_chan_dep_data_7;
    wire [32:0] token_out_vec_7;
    wire dl_detect_out_7;
    wire dep_chan_vld_0_7;
    wire [39:0] dep_chan_data_0_7;
    wire token_0_7;
    wire dep_chan_vld_1_7;
    wire [39:0] dep_chan_data_1_7;
    wire token_1_7;
    wire dep_chan_vld_3_7;
    wire [39:0] dep_chan_data_3_7;
    wire token_3_7;
    wire dep_chan_vld_6_7;
    wire [39:0] dep_chan_data_6_7;
    wire token_6_7;
    wire dep_chan_vld_8_7;
    wire [39:0] dep_chan_data_8_7;
    wire token_8_7;
    wire dep_chan_vld_9_7;
    wire [39:0] dep_chan_data_9_7;
    wire token_9_7;
    wire dep_chan_vld_10_7;
    wire [39:0] dep_chan_data_10_7;
    wire token_10_7;
    wire dep_chan_vld_11_7;
    wire [39:0] dep_chan_data_11_7;
    wire token_11_7;
    wire dep_chan_vld_12_7;
    wire [39:0] dep_chan_data_12_7;
    wire token_12_7;
    wire dep_chan_vld_13_7;
    wire [39:0] dep_chan_data_13_7;
    wire token_13_7;
    wire dep_chan_vld_14_7;
    wire [39:0] dep_chan_data_14_7;
    wire token_14_7;
    wire dep_chan_vld_15_7;
    wire [39:0] dep_chan_data_15_7;
    wire token_15_7;
    wire dep_chan_vld_16_7;
    wire [39:0] dep_chan_data_16_7;
    wire token_16_7;
    wire dep_chan_vld_17_7;
    wire [39:0] dep_chan_data_17_7;
    wire token_17_7;
    wire dep_chan_vld_18_7;
    wire [39:0] dep_chan_data_18_7;
    wire token_18_7;
    wire dep_chan_vld_19_7;
    wire [39:0] dep_chan_data_19_7;
    wire token_19_7;
    wire dep_chan_vld_20_7;
    wire [39:0] dep_chan_data_20_7;
    wire token_20_7;
    wire dep_chan_vld_21_7;
    wire [39:0] dep_chan_data_21_7;
    wire token_21_7;
    wire dep_chan_vld_22_7;
    wire [39:0] dep_chan_data_22_7;
    wire token_22_7;
    wire dep_chan_vld_23_7;
    wire [39:0] dep_chan_data_23_7;
    wire token_23_7;
    wire dep_chan_vld_24_7;
    wire [39:0] dep_chan_data_24_7;
    wire token_24_7;
    wire dep_chan_vld_25_7;
    wire [39:0] dep_chan_data_25_7;
    wire token_25_7;
    wire dep_chan_vld_26_7;
    wire [39:0] dep_chan_data_26_7;
    wire token_26_7;
    wire dep_chan_vld_27_7;
    wire [39:0] dep_chan_data_27_7;
    wire token_27_7;
    wire dep_chan_vld_28_7;
    wire [39:0] dep_chan_data_28_7;
    wire token_28_7;
    wire dep_chan_vld_29_7;
    wire [39:0] dep_chan_data_29_7;
    wire token_29_7;
    wire dep_chan_vld_30_7;
    wire [39:0] dep_chan_data_30_7;
    wire token_30_7;
    wire dep_chan_vld_31_7;
    wire [39:0] dep_chan_data_31_7;
    wire token_31_7;
    wire dep_chan_vld_32_7;
    wire [39:0] dep_chan_data_32_7;
    wire token_32_7;
    wire dep_chan_vld_33_7;
    wire [39:0] dep_chan_data_33_7;
    wire token_33_7;
    wire dep_chan_vld_34_7;
    wire [39:0] dep_chan_data_34_7;
    wire token_34_7;
    wire dep_chan_vld_35_7;
    wire [39:0] dep_chan_data_35_7;
    wire token_35_7;
    wire dep_chan_vld_36_7;
    wire [39:0] dep_chan_data_36_7;
    wire token_36_7;
    wire [32:0] proc_8_data_FIFO_blk;
    wire [32:0] proc_8_data_PIPO_blk;
    wire [32:0] proc_8_start_FIFO_blk;
    wire [32:0] proc_8_TLF_FIFO_blk;
    wire [32:0] proc_8_input_sync_blk;
    wire [32:0] proc_8_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_8;
    reg [32:0] proc_dep_vld_vec_8_reg;
    wire [32:0] in_chan_dep_vld_vec_8;
    wire [1319:0] in_chan_dep_data_vec_8;
    wire [32:0] token_in_vec_8;
    wire [32:0] out_chan_dep_vld_vec_8;
    wire [39:0] out_chan_dep_data_8;
    wire [32:0] token_out_vec_8;
    wire dl_detect_out_8;
    wire dep_chan_vld_0_8;
    wire [39:0] dep_chan_data_0_8;
    wire token_0_8;
    wire dep_chan_vld_1_8;
    wire [39:0] dep_chan_data_1_8;
    wire token_1_8;
    wire dep_chan_vld_3_8;
    wire [39:0] dep_chan_data_3_8;
    wire token_3_8;
    wire dep_chan_vld_6_8;
    wire [39:0] dep_chan_data_6_8;
    wire token_6_8;
    wire dep_chan_vld_7_8;
    wire [39:0] dep_chan_data_7_8;
    wire token_7_8;
    wire dep_chan_vld_9_8;
    wire [39:0] dep_chan_data_9_8;
    wire token_9_8;
    wire dep_chan_vld_10_8;
    wire [39:0] dep_chan_data_10_8;
    wire token_10_8;
    wire dep_chan_vld_11_8;
    wire [39:0] dep_chan_data_11_8;
    wire token_11_8;
    wire dep_chan_vld_12_8;
    wire [39:0] dep_chan_data_12_8;
    wire token_12_8;
    wire dep_chan_vld_13_8;
    wire [39:0] dep_chan_data_13_8;
    wire token_13_8;
    wire dep_chan_vld_14_8;
    wire [39:0] dep_chan_data_14_8;
    wire token_14_8;
    wire dep_chan_vld_15_8;
    wire [39:0] dep_chan_data_15_8;
    wire token_15_8;
    wire dep_chan_vld_16_8;
    wire [39:0] dep_chan_data_16_8;
    wire token_16_8;
    wire dep_chan_vld_17_8;
    wire [39:0] dep_chan_data_17_8;
    wire token_17_8;
    wire dep_chan_vld_18_8;
    wire [39:0] dep_chan_data_18_8;
    wire token_18_8;
    wire dep_chan_vld_19_8;
    wire [39:0] dep_chan_data_19_8;
    wire token_19_8;
    wire dep_chan_vld_20_8;
    wire [39:0] dep_chan_data_20_8;
    wire token_20_8;
    wire dep_chan_vld_21_8;
    wire [39:0] dep_chan_data_21_8;
    wire token_21_8;
    wire dep_chan_vld_22_8;
    wire [39:0] dep_chan_data_22_8;
    wire token_22_8;
    wire dep_chan_vld_23_8;
    wire [39:0] dep_chan_data_23_8;
    wire token_23_8;
    wire dep_chan_vld_24_8;
    wire [39:0] dep_chan_data_24_8;
    wire token_24_8;
    wire dep_chan_vld_25_8;
    wire [39:0] dep_chan_data_25_8;
    wire token_25_8;
    wire dep_chan_vld_26_8;
    wire [39:0] dep_chan_data_26_8;
    wire token_26_8;
    wire dep_chan_vld_27_8;
    wire [39:0] dep_chan_data_27_8;
    wire token_27_8;
    wire dep_chan_vld_28_8;
    wire [39:0] dep_chan_data_28_8;
    wire token_28_8;
    wire dep_chan_vld_29_8;
    wire [39:0] dep_chan_data_29_8;
    wire token_29_8;
    wire dep_chan_vld_30_8;
    wire [39:0] dep_chan_data_30_8;
    wire token_30_8;
    wire dep_chan_vld_31_8;
    wire [39:0] dep_chan_data_31_8;
    wire token_31_8;
    wire dep_chan_vld_32_8;
    wire [39:0] dep_chan_data_32_8;
    wire token_32_8;
    wire dep_chan_vld_33_8;
    wire [39:0] dep_chan_data_33_8;
    wire token_33_8;
    wire dep_chan_vld_34_8;
    wire [39:0] dep_chan_data_34_8;
    wire token_34_8;
    wire dep_chan_vld_35_8;
    wire [39:0] dep_chan_data_35_8;
    wire token_35_8;
    wire dep_chan_vld_36_8;
    wire [39:0] dep_chan_data_36_8;
    wire token_36_8;
    wire [32:0] proc_9_data_FIFO_blk;
    wire [32:0] proc_9_data_PIPO_blk;
    wire [32:0] proc_9_start_FIFO_blk;
    wire [32:0] proc_9_TLF_FIFO_blk;
    wire [32:0] proc_9_input_sync_blk;
    wire [32:0] proc_9_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_9;
    reg [32:0] proc_dep_vld_vec_9_reg;
    wire [32:0] in_chan_dep_vld_vec_9;
    wire [1319:0] in_chan_dep_data_vec_9;
    wire [32:0] token_in_vec_9;
    wire [32:0] out_chan_dep_vld_vec_9;
    wire [39:0] out_chan_dep_data_9;
    wire [32:0] token_out_vec_9;
    wire dl_detect_out_9;
    wire dep_chan_vld_0_9;
    wire [39:0] dep_chan_data_0_9;
    wire token_0_9;
    wire dep_chan_vld_1_9;
    wire [39:0] dep_chan_data_1_9;
    wire token_1_9;
    wire dep_chan_vld_3_9;
    wire [39:0] dep_chan_data_3_9;
    wire token_3_9;
    wire dep_chan_vld_6_9;
    wire [39:0] dep_chan_data_6_9;
    wire token_6_9;
    wire dep_chan_vld_7_9;
    wire [39:0] dep_chan_data_7_9;
    wire token_7_9;
    wire dep_chan_vld_8_9;
    wire [39:0] dep_chan_data_8_9;
    wire token_8_9;
    wire dep_chan_vld_10_9;
    wire [39:0] dep_chan_data_10_9;
    wire token_10_9;
    wire dep_chan_vld_11_9;
    wire [39:0] dep_chan_data_11_9;
    wire token_11_9;
    wire dep_chan_vld_12_9;
    wire [39:0] dep_chan_data_12_9;
    wire token_12_9;
    wire dep_chan_vld_13_9;
    wire [39:0] dep_chan_data_13_9;
    wire token_13_9;
    wire dep_chan_vld_14_9;
    wire [39:0] dep_chan_data_14_9;
    wire token_14_9;
    wire dep_chan_vld_15_9;
    wire [39:0] dep_chan_data_15_9;
    wire token_15_9;
    wire dep_chan_vld_16_9;
    wire [39:0] dep_chan_data_16_9;
    wire token_16_9;
    wire dep_chan_vld_17_9;
    wire [39:0] dep_chan_data_17_9;
    wire token_17_9;
    wire dep_chan_vld_18_9;
    wire [39:0] dep_chan_data_18_9;
    wire token_18_9;
    wire dep_chan_vld_19_9;
    wire [39:0] dep_chan_data_19_9;
    wire token_19_9;
    wire dep_chan_vld_20_9;
    wire [39:0] dep_chan_data_20_9;
    wire token_20_9;
    wire dep_chan_vld_21_9;
    wire [39:0] dep_chan_data_21_9;
    wire token_21_9;
    wire dep_chan_vld_22_9;
    wire [39:0] dep_chan_data_22_9;
    wire token_22_9;
    wire dep_chan_vld_23_9;
    wire [39:0] dep_chan_data_23_9;
    wire token_23_9;
    wire dep_chan_vld_24_9;
    wire [39:0] dep_chan_data_24_9;
    wire token_24_9;
    wire dep_chan_vld_25_9;
    wire [39:0] dep_chan_data_25_9;
    wire token_25_9;
    wire dep_chan_vld_26_9;
    wire [39:0] dep_chan_data_26_9;
    wire token_26_9;
    wire dep_chan_vld_27_9;
    wire [39:0] dep_chan_data_27_9;
    wire token_27_9;
    wire dep_chan_vld_28_9;
    wire [39:0] dep_chan_data_28_9;
    wire token_28_9;
    wire dep_chan_vld_29_9;
    wire [39:0] dep_chan_data_29_9;
    wire token_29_9;
    wire dep_chan_vld_30_9;
    wire [39:0] dep_chan_data_30_9;
    wire token_30_9;
    wire dep_chan_vld_31_9;
    wire [39:0] dep_chan_data_31_9;
    wire token_31_9;
    wire dep_chan_vld_32_9;
    wire [39:0] dep_chan_data_32_9;
    wire token_32_9;
    wire dep_chan_vld_33_9;
    wire [39:0] dep_chan_data_33_9;
    wire token_33_9;
    wire dep_chan_vld_34_9;
    wire [39:0] dep_chan_data_34_9;
    wire token_34_9;
    wire dep_chan_vld_35_9;
    wire [39:0] dep_chan_data_35_9;
    wire token_35_9;
    wire dep_chan_vld_36_9;
    wire [39:0] dep_chan_data_36_9;
    wire token_36_9;
    wire [32:0] proc_10_data_FIFO_blk;
    wire [32:0] proc_10_data_PIPO_blk;
    wire [32:0] proc_10_start_FIFO_blk;
    wire [32:0] proc_10_TLF_FIFO_blk;
    wire [32:0] proc_10_input_sync_blk;
    wire [32:0] proc_10_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_10;
    reg [32:0] proc_dep_vld_vec_10_reg;
    wire [32:0] in_chan_dep_vld_vec_10;
    wire [1319:0] in_chan_dep_data_vec_10;
    wire [32:0] token_in_vec_10;
    wire [32:0] out_chan_dep_vld_vec_10;
    wire [39:0] out_chan_dep_data_10;
    wire [32:0] token_out_vec_10;
    wire dl_detect_out_10;
    wire dep_chan_vld_0_10;
    wire [39:0] dep_chan_data_0_10;
    wire token_0_10;
    wire dep_chan_vld_1_10;
    wire [39:0] dep_chan_data_1_10;
    wire token_1_10;
    wire dep_chan_vld_3_10;
    wire [39:0] dep_chan_data_3_10;
    wire token_3_10;
    wire dep_chan_vld_6_10;
    wire [39:0] dep_chan_data_6_10;
    wire token_6_10;
    wire dep_chan_vld_7_10;
    wire [39:0] dep_chan_data_7_10;
    wire token_7_10;
    wire dep_chan_vld_8_10;
    wire [39:0] dep_chan_data_8_10;
    wire token_8_10;
    wire dep_chan_vld_9_10;
    wire [39:0] dep_chan_data_9_10;
    wire token_9_10;
    wire dep_chan_vld_11_10;
    wire [39:0] dep_chan_data_11_10;
    wire token_11_10;
    wire dep_chan_vld_12_10;
    wire [39:0] dep_chan_data_12_10;
    wire token_12_10;
    wire dep_chan_vld_13_10;
    wire [39:0] dep_chan_data_13_10;
    wire token_13_10;
    wire dep_chan_vld_14_10;
    wire [39:0] dep_chan_data_14_10;
    wire token_14_10;
    wire dep_chan_vld_15_10;
    wire [39:0] dep_chan_data_15_10;
    wire token_15_10;
    wire dep_chan_vld_16_10;
    wire [39:0] dep_chan_data_16_10;
    wire token_16_10;
    wire dep_chan_vld_17_10;
    wire [39:0] dep_chan_data_17_10;
    wire token_17_10;
    wire dep_chan_vld_18_10;
    wire [39:0] dep_chan_data_18_10;
    wire token_18_10;
    wire dep_chan_vld_19_10;
    wire [39:0] dep_chan_data_19_10;
    wire token_19_10;
    wire dep_chan_vld_20_10;
    wire [39:0] dep_chan_data_20_10;
    wire token_20_10;
    wire dep_chan_vld_21_10;
    wire [39:0] dep_chan_data_21_10;
    wire token_21_10;
    wire dep_chan_vld_22_10;
    wire [39:0] dep_chan_data_22_10;
    wire token_22_10;
    wire dep_chan_vld_23_10;
    wire [39:0] dep_chan_data_23_10;
    wire token_23_10;
    wire dep_chan_vld_24_10;
    wire [39:0] dep_chan_data_24_10;
    wire token_24_10;
    wire dep_chan_vld_25_10;
    wire [39:0] dep_chan_data_25_10;
    wire token_25_10;
    wire dep_chan_vld_26_10;
    wire [39:0] dep_chan_data_26_10;
    wire token_26_10;
    wire dep_chan_vld_27_10;
    wire [39:0] dep_chan_data_27_10;
    wire token_27_10;
    wire dep_chan_vld_28_10;
    wire [39:0] dep_chan_data_28_10;
    wire token_28_10;
    wire dep_chan_vld_29_10;
    wire [39:0] dep_chan_data_29_10;
    wire token_29_10;
    wire dep_chan_vld_30_10;
    wire [39:0] dep_chan_data_30_10;
    wire token_30_10;
    wire dep_chan_vld_31_10;
    wire [39:0] dep_chan_data_31_10;
    wire token_31_10;
    wire dep_chan_vld_32_10;
    wire [39:0] dep_chan_data_32_10;
    wire token_32_10;
    wire dep_chan_vld_33_10;
    wire [39:0] dep_chan_data_33_10;
    wire token_33_10;
    wire dep_chan_vld_34_10;
    wire [39:0] dep_chan_data_34_10;
    wire token_34_10;
    wire dep_chan_vld_35_10;
    wire [39:0] dep_chan_data_35_10;
    wire token_35_10;
    wire dep_chan_vld_36_10;
    wire [39:0] dep_chan_data_36_10;
    wire token_36_10;
    wire [32:0] proc_11_data_FIFO_blk;
    wire [32:0] proc_11_data_PIPO_blk;
    wire [32:0] proc_11_start_FIFO_blk;
    wire [32:0] proc_11_TLF_FIFO_blk;
    wire [32:0] proc_11_input_sync_blk;
    wire [32:0] proc_11_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_11;
    reg [32:0] proc_dep_vld_vec_11_reg;
    wire [32:0] in_chan_dep_vld_vec_11;
    wire [1319:0] in_chan_dep_data_vec_11;
    wire [32:0] token_in_vec_11;
    wire [32:0] out_chan_dep_vld_vec_11;
    wire [39:0] out_chan_dep_data_11;
    wire [32:0] token_out_vec_11;
    wire dl_detect_out_11;
    wire dep_chan_vld_0_11;
    wire [39:0] dep_chan_data_0_11;
    wire token_0_11;
    wire dep_chan_vld_1_11;
    wire [39:0] dep_chan_data_1_11;
    wire token_1_11;
    wire dep_chan_vld_3_11;
    wire [39:0] dep_chan_data_3_11;
    wire token_3_11;
    wire dep_chan_vld_6_11;
    wire [39:0] dep_chan_data_6_11;
    wire token_6_11;
    wire dep_chan_vld_7_11;
    wire [39:0] dep_chan_data_7_11;
    wire token_7_11;
    wire dep_chan_vld_8_11;
    wire [39:0] dep_chan_data_8_11;
    wire token_8_11;
    wire dep_chan_vld_9_11;
    wire [39:0] dep_chan_data_9_11;
    wire token_9_11;
    wire dep_chan_vld_10_11;
    wire [39:0] dep_chan_data_10_11;
    wire token_10_11;
    wire dep_chan_vld_12_11;
    wire [39:0] dep_chan_data_12_11;
    wire token_12_11;
    wire dep_chan_vld_13_11;
    wire [39:0] dep_chan_data_13_11;
    wire token_13_11;
    wire dep_chan_vld_14_11;
    wire [39:0] dep_chan_data_14_11;
    wire token_14_11;
    wire dep_chan_vld_15_11;
    wire [39:0] dep_chan_data_15_11;
    wire token_15_11;
    wire dep_chan_vld_16_11;
    wire [39:0] dep_chan_data_16_11;
    wire token_16_11;
    wire dep_chan_vld_17_11;
    wire [39:0] dep_chan_data_17_11;
    wire token_17_11;
    wire dep_chan_vld_18_11;
    wire [39:0] dep_chan_data_18_11;
    wire token_18_11;
    wire dep_chan_vld_19_11;
    wire [39:0] dep_chan_data_19_11;
    wire token_19_11;
    wire dep_chan_vld_20_11;
    wire [39:0] dep_chan_data_20_11;
    wire token_20_11;
    wire dep_chan_vld_21_11;
    wire [39:0] dep_chan_data_21_11;
    wire token_21_11;
    wire dep_chan_vld_22_11;
    wire [39:0] dep_chan_data_22_11;
    wire token_22_11;
    wire dep_chan_vld_23_11;
    wire [39:0] dep_chan_data_23_11;
    wire token_23_11;
    wire dep_chan_vld_24_11;
    wire [39:0] dep_chan_data_24_11;
    wire token_24_11;
    wire dep_chan_vld_25_11;
    wire [39:0] dep_chan_data_25_11;
    wire token_25_11;
    wire dep_chan_vld_26_11;
    wire [39:0] dep_chan_data_26_11;
    wire token_26_11;
    wire dep_chan_vld_27_11;
    wire [39:0] dep_chan_data_27_11;
    wire token_27_11;
    wire dep_chan_vld_28_11;
    wire [39:0] dep_chan_data_28_11;
    wire token_28_11;
    wire dep_chan_vld_29_11;
    wire [39:0] dep_chan_data_29_11;
    wire token_29_11;
    wire dep_chan_vld_30_11;
    wire [39:0] dep_chan_data_30_11;
    wire token_30_11;
    wire dep_chan_vld_31_11;
    wire [39:0] dep_chan_data_31_11;
    wire token_31_11;
    wire dep_chan_vld_32_11;
    wire [39:0] dep_chan_data_32_11;
    wire token_32_11;
    wire dep_chan_vld_33_11;
    wire [39:0] dep_chan_data_33_11;
    wire token_33_11;
    wire dep_chan_vld_34_11;
    wire [39:0] dep_chan_data_34_11;
    wire token_34_11;
    wire dep_chan_vld_35_11;
    wire [39:0] dep_chan_data_35_11;
    wire token_35_11;
    wire dep_chan_vld_36_11;
    wire [39:0] dep_chan_data_36_11;
    wire token_36_11;
    wire [32:0] proc_12_data_FIFO_blk;
    wire [32:0] proc_12_data_PIPO_blk;
    wire [32:0] proc_12_start_FIFO_blk;
    wire [32:0] proc_12_TLF_FIFO_blk;
    wire [32:0] proc_12_input_sync_blk;
    wire [32:0] proc_12_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_12;
    reg [32:0] proc_dep_vld_vec_12_reg;
    wire [32:0] in_chan_dep_vld_vec_12;
    wire [1319:0] in_chan_dep_data_vec_12;
    wire [32:0] token_in_vec_12;
    wire [32:0] out_chan_dep_vld_vec_12;
    wire [39:0] out_chan_dep_data_12;
    wire [32:0] token_out_vec_12;
    wire dl_detect_out_12;
    wire dep_chan_vld_0_12;
    wire [39:0] dep_chan_data_0_12;
    wire token_0_12;
    wire dep_chan_vld_1_12;
    wire [39:0] dep_chan_data_1_12;
    wire token_1_12;
    wire dep_chan_vld_3_12;
    wire [39:0] dep_chan_data_3_12;
    wire token_3_12;
    wire dep_chan_vld_6_12;
    wire [39:0] dep_chan_data_6_12;
    wire token_6_12;
    wire dep_chan_vld_7_12;
    wire [39:0] dep_chan_data_7_12;
    wire token_7_12;
    wire dep_chan_vld_8_12;
    wire [39:0] dep_chan_data_8_12;
    wire token_8_12;
    wire dep_chan_vld_9_12;
    wire [39:0] dep_chan_data_9_12;
    wire token_9_12;
    wire dep_chan_vld_10_12;
    wire [39:0] dep_chan_data_10_12;
    wire token_10_12;
    wire dep_chan_vld_11_12;
    wire [39:0] dep_chan_data_11_12;
    wire token_11_12;
    wire dep_chan_vld_13_12;
    wire [39:0] dep_chan_data_13_12;
    wire token_13_12;
    wire dep_chan_vld_14_12;
    wire [39:0] dep_chan_data_14_12;
    wire token_14_12;
    wire dep_chan_vld_15_12;
    wire [39:0] dep_chan_data_15_12;
    wire token_15_12;
    wire dep_chan_vld_16_12;
    wire [39:0] dep_chan_data_16_12;
    wire token_16_12;
    wire dep_chan_vld_17_12;
    wire [39:0] dep_chan_data_17_12;
    wire token_17_12;
    wire dep_chan_vld_18_12;
    wire [39:0] dep_chan_data_18_12;
    wire token_18_12;
    wire dep_chan_vld_19_12;
    wire [39:0] dep_chan_data_19_12;
    wire token_19_12;
    wire dep_chan_vld_20_12;
    wire [39:0] dep_chan_data_20_12;
    wire token_20_12;
    wire dep_chan_vld_21_12;
    wire [39:0] dep_chan_data_21_12;
    wire token_21_12;
    wire dep_chan_vld_22_12;
    wire [39:0] dep_chan_data_22_12;
    wire token_22_12;
    wire dep_chan_vld_23_12;
    wire [39:0] dep_chan_data_23_12;
    wire token_23_12;
    wire dep_chan_vld_24_12;
    wire [39:0] dep_chan_data_24_12;
    wire token_24_12;
    wire dep_chan_vld_25_12;
    wire [39:0] dep_chan_data_25_12;
    wire token_25_12;
    wire dep_chan_vld_26_12;
    wire [39:0] dep_chan_data_26_12;
    wire token_26_12;
    wire dep_chan_vld_27_12;
    wire [39:0] dep_chan_data_27_12;
    wire token_27_12;
    wire dep_chan_vld_28_12;
    wire [39:0] dep_chan_data_28_12;
    wire token_28_12;
    wire dep_chan_vld_29_12;
    wire [39:0] dep_chan_data_29_12;
    wire token_29_12;
    wire dep_chan_vld_30_12;
    wire [39:0] dep_chan_data_30_12;
    wire token_30_12;
    wire dep_chan_vld_31_12;
    wire [39:0] dep_chan_data_31_12;
    wire token_31_12;
    wire dep_chan_vld_32_12;
    wire [39:0] dep_chan_data_32_12;
    wire token_32_12;
    wire dep_chan_vld_33_12;
    wire [39:0] dep_chan_data_33_12;
    wire token_33_12;
    wire dep_chan_vld_34_12;
    wire [39:0] dep_chan_data_34_12;
    wire token_34_12;
    wire dep_chan_vld_35_12;
    wire [39:0] dep_chan_data_35_12;
    wire token_35_12;
    wire dep_chan_vld_36_12;
    wire [39:0] dep_chan_data_36_12;
    wire token_36_12;
    wire [32:0] proc_13_data_FIFO_blk;
    wire [32:0] proc_13_data_PIPO_blk;
    wire [32:0] proc_13_start_FIFO_blk;
    wire [32:0] proc_13_TLF_FIFO_blk;
    wire [32:0] proc_13_input_sync_blk;
    wire [32:0] proc_13_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_13;
    reg [32:0] proc_dep_vld_vec_13_reg;
    wire [32:0] in_chan_dep_vld_vec_13;
    wire [1319:0] in_chan_dep_data_vec_13;
    wire [32:0] token_in_vec_13;
    wire [32:0] out_chan_dep_vld_vec_13;
    wire [39:0] out_chan_dep_data_13;
    wire [32:0] token_out_vec_13;
    wire dl_detect_out_13;
    wire dep_chan_vld_0_13;
    wire [39:0] dep_chan_data_0_13;
    wire token_0_13;
    wire dep_chan_vld_1_13;
    wire [39:0] dep_chan_data_1_13;
    wire token_1_13;
    wire dep_chan_vld_3_13;
    wire [39:0] dep_chan_data_3_13;
    wire token_3_13;
    wire dep_chan_vld_6_13;
    wire [39:0] dep_chan_data_6_13;
    wire token_6_13;
    wire dep_chan_vld_7_13;
    wire [39:0] dep_chan_data_7_13;
    wire token_7_13;
    wire dep_chan_vld_8_13;
    wire [39:0] dep_chan_data_8_13;
    wire token_8_13;
    wire dep_chan_vld_9_13;
    wire [39:0] dep_chan_data_9_13;
    wire token_9_13;
    wire dep_chan_vld_10_13;
    wire [39:0] dep_chan_data_10_13;
    wire token_10_13;
    wire dep_chan_vld_11_13;
    wire [39:0] dep_chan_data_11_13;
    wire token_11_13;
    wire dep_chan_vld_12_13;
    wire [39:0] dep_chan_data_12_13;
    wire token_12_13;
    wire dep_chan_vld_14_13;
    wire [39:0] dep_chan_data_14_13;
    wire token_14_13;
    wire dep_chan_vld_15_13;
    wire [39:0] dep_chan_data_15_13;
    wire token_15_13;
    wire dep_chan_vld_16_13;
    wire [39:0] dep_chan_data_16_13;
    wire token_16_13;
    wire dep_chan_vld_17_13;
    wire [39:0] dep_chan_data_17_13;
    wire token_17_13;
    wire dep_chan_vld_18_13;
    wire [39:0] dep_chan_data_18_13;
    wire token_18_13;
    wire dep_chan_vld_19_13;
    wire [39:0] dep_chan_data_19_13;
    wire token_19_13;
    wire dep_chan_vld_20_13;
    wire [39:0] dep_chan_data_20_13;
    wire token_20_13;
    wire dep_chan_vld_21_13;
    wire [39:0] dep_chan_data_21_13;
    wire token_21_13;
    wire dep_chan_vld_22_13;
    wire [39:0] dep_chan_data_22_13;
    wire token_22_13;
    wire dep_chan_vld_23_13;
    wire [39:0] dep_chan_data_23_13;
    wire token_23_13;
    wire dep_chan_vld_24_13;
    wire [39:0] dep_chan_data_24_13;
    wire token_24_13;
    wire dep_chan_vld_25_13;
    wire [39:0] dep_chan_data_25_13;
    wire token_25_13;
    wire dep_chan_vld_26_13;
    wire [39:0] dep_chan_data_26_13;
    wire token_26_13;
    wire dep_chan_vld_27_13;
    wire [39:0] dep_chan_data_27_13;
    wire token_27_13;
    wire dep_chan_vld_28_13;
    wire [39:0] dep_chan_data_28_13;
    wire token_28_13;
    wire dep_chan_vld_29_13;
    wire [39:0] dep_chan_data_29_13;
    wire token_29_13;
    wire dep_chan_vld_30_13;
    wire [39:0] dep_chan_data_30_13;
    wire token_30_13;
    wire dep_chan_vld_31_13;
    wire [39:0] dep_chan_data_31_13;
    wire token_31_13;
    wire dep_chan_vld_32_13;
    wire [39:0] dep_chan_data_32_13;
    wire token_32_13;
    wire dep_chan_vld_33_13;
    wire [39:0] dep_chan_data_33_13;
    wire token_33_13;
    wire dep_chan_vld_34_13;
    wire [39:0] dep_chan_data_34_13;
    wire token_34_13;
    wire dep_chan_vld_35_13;
    wire [39:0] dep_chan_data_35_13;
    wire token_35_13;
    wire dep_chan_vld_36_13;
    wire [39:0] dep_chan_data_36_13;
    wire token_36_13;
    wire [32:0] proc_14_data_FIFO_blk;
    wire [32:0] proc_14_data_PIPO_blk;
    wire [32:0] proc_14_start_FIFO_blk;
    wire [32:0] proc_14_TLF_FIFO_blk;
    wire [32:0] proc_14_input_sync_blk;
    wire [32:0] proc_14_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_14;
    reg [32:0] proc_dep_vld_vec_14_reg;
    wire [32:0] in_chan_dep_vld_vec_14;
    wire [1319:0] in_chan_dep_data_vec_14;
    wire [32:0] token_in_vec_14;
    wire [32:0] out_chan_dep_vld_vec_14;
    wire [39:0] out_chan_dep_data_14;
    wire [32:0] token_out_vec_14;
    wire dl_detect_out_14;
    wire dep_chan_vld_0_14;
    wire [39:0] dep_chan_data_0_14;
    wire token_0_14;
    wire dep_chan_vld_1_14;
    wire [39:0] dep_chan_data_1_14;
    wire token_1_14;
    wire dep_chan_vld_3_14;
    wire [39:0] dep_chan_data_3_14;
    wire token_3_14;
    wire dep_chan_vld_6_14;
    wire [39:0] dep_chan_data_6_14;
    wire token_6_14;
    wire dep_chan_vld_7_14;
    wire [39:0] dep_chan_data_7_14;
    wire token_7_14;
    wire dep_chan_vld_8_14;
    wire [39:0] dep_chan_data_8_14;
    wire token_8_14;
    wire dep_chan_vld_9_14;
    wire [39:0] dep_chan_data_9_14;
    wire token_9_14;
    wire dep_chan_vld_10_14;
    wire [39:0] dep_chan_data_10_14;
    wire token_10_14;
    wire dep_chan_vld_11_14;
    wire [39:0] dep_chan_data_11_14;
    wire token_11_14;
    wire dep_chan_vld_12_14;
    wire [39:0] dep_chan_data_12_14;
    wire token_12_14;
    wire dep_chan_vld_13_14;
    wire [39:0] dep_chan_data_13_14;
    wire token_13_14;
    wire dep_chan_vld_15_14;
    wire [39:0] dep_chan_data_15_14;
    wire token_15_14;
    wire dep_chan_vld_16_14;
    wire [39:0] dep_chan_data_16_14;
    wire token_16_14;
    wire dep_chan_vld_17_14;
    wire [39:0] dep_chan_data_17_14;
    wire token_17_14;
    wire dep_chan_vld_18_14;
    wire [39:0] dep_chan_data_18_14;
    wire token_18_14;
    wire dep_chan_vld_19_14;
    wire [39:0] dep_chan_data_19_14;
    wire token_19_14;
    wire dep_chan_vld_20_14;
    wire [39:0] dep_chan_data_20_14;
    wire token_20_14;
    wire dep_chan_vld_21_14;
    wire [39:0] dep_chan_data_21_14;
    wire token_21_14;
    wire dep_chan_vld_22_14;
    wire [39:0] dep_chan_data_22_14;
    wire token_22_14;
    wire dep_chan_vld_23_14;
    wire [39:0] dep_chan_data_23_14;
    wire token_23_14;
    wire dep_chan_vld_24_14;
    wire [39:0] dep_chan_data_24_14;
    wire token_24_14;
    wire dep_chan_vld_25_14;
    wire [39:0] dep_chan_data_25_14;
    wire token_25_14;
    wire dep_chan_vld_26_14;
    wire [39:0] dep_chan_data_26_14;
    wire token_26_14;
    wire dep_chan_vld_27_14;
    wire [39:0] dep_chan_data_27_14;
    wire token_27_14;
    wire dep_chan_vld_28_14;
    wire [39:0] dep_chan_data_28_14;
    wire token_28_14;
    wire dep_chan_vld_29_14;
    wire [39:0] dep_chan_data_29_14;
    wire token_29_14;
    wire dep_chan_vld_30_14;
    wire [39:0] dep_chan_data_30_14;
    wire token_30_14;
    wire dep_chan_vld_31_14;
    wire [39:0] dep_chan_data_31_14;
    wire token_31_14;
    wire dep_chan_vld_32_14;
    wire [39:0] dep_chan_data_32_14;
    wire token_32_14;
    wire dep_chan_vld_33_14;
    wire [39:0] dep_chan_data_33_14;
    wire token_33_14;
    wire dep_chan_vld_34_14;
    wire [39:0] dep_chan_data_34_14;
    wire token_34_14;
    wire dep_chan_vld_35_14;
    wire [39:0] dep_chan_data_35_14;
    wire token_35_14;
    wire dep_chan_vld_36_14;
    wire [39:0] dep_chan_data_36_14;
    wire token_36_14;
    wire [32:0] proc_15_data_FIFO_blk;
    wire [32:0] proc_15_data_PIPO_blk;
    wire [32:0] proc_15_start_FIFO_blk;
    wire [32:0] proc_15_TLF_FIFO_blk;
    wire [32:0] proc_15_input_sync_blk;
    wire [32:0] proc_15_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_15;
    reg [32:0] proc_dep_vld_vec_15_reg;
    wire [32:0] in_chan_dep_vld_vec_15;
    wire [1319:0] in_chan_dep_data_vec_15;
    wire [32:0] token_in_vec_15;
    wire [32:0] out_chan_dep_vld_vec_15;
    wire [39:0] out_chan_dep_data_15;
    wire [32:0] token_out_vec_15;
    wire dl_detect_out_15;
    wire dep_chan_vld_0_15;
    wire [39:0] dep_chan_data_0_15;
    wire token_0_15;
    wire dep_chan_vld_1_15;
    wire [39:0] dep_chan_data_1_15;
    wire token_1_15;
    wire dep_chan_vld_3_15;
    wire [39:0] dep_chan_data_3_15;
    wire token_3_15;
    wire dep_chan_vld_6_15;
    wire [39:0] dep_chan_data_6_15;
    wire token_6_15;
    wire dep_chan_vld_7_15;
    wire [39:0] dep_chan_data_7_15;
    wire token_7_15;
    wire dep_chan_vld_8_15;
    wire [39:0] dep_chan_data_8_15;
    wire token_8_15;
    wire dep_chan_vld_9_15;
    wire [39:0] dep_chan_data_9_15;
    wire token_9_15;
    wire dep_chan_vld_10_15;
    wire [39:0] dep_chan_data_10_15;
    wire token_10_15;
    wire dep_chan_vld_11_15;
    wire [39:0] dep_chan_data_11_15;
    wire token_11_15;
    wire dep_chan_vld_12_15;
    wire [39:0] dep_chan_data_12_15;
    wire token_12_15;
    wire dep_chan_vld_13_15;
    wire [39:0] dep_chan_data_13_15;
    wire token_13_15;
    wire dep_chan_vld_14_15;
    wire [39:0] dep_chan_data_14_15;
    wire token_14_15;
    wire dep_chan_vld_16_15;
    wire [39:0] dep_chan_data_16_15;
    wire token_16_15;
    wire dep_chan_vld_17_15;
    wire [39:0] dep_chan_data_17_15;
    wire token_17_15;
    wire dep_chan_vld_18_15;
    wire [39:0] dep_chan_data_18_15;
    wire token_18_15;
    wire dep_chan_vld_19_15;
    wire [39:0] dep_chan_data_19_15;
    wire token_19_15;
    wire dep_chan_vld_20_15;
    wire [39:0] dep_chan_data_20_15;
    wire token_20_15;
    wire dep_chan_vld_21_15;
    wire [39:0] dep_chan_data_21_15;
    wire token_21_15;
    wire dep_chan_vld_22_15;
    wire [39:0] dep_chan_data_22_15;
    wire token_22_15;
    wire dep_chan_vld_23_15;
    wire [39:0] dep_chan_data_23_15;
    wire token_23_15;
    wire dep_chan_vld_24_15;
    wire [39:0] dep_chan_data_24_15;
    wire token_24_15;
    wire dep_chan_vld_25_15;
    wire [39:0] dep_chan_data_25_15;
    wire token_25_15;
    wire dep_chan_vld_26_15;
    wire [39:0] dep_chan_data_26_15;
    wire token_26_15;
    wire dep_chan_vld_27_15;
    wire [39:0] dep_chan_data_27_15;
    wire token_27_15;
    wire dep_chan_vld_28_15;
    wire [39:0] dep_chan_data_28_15;
    wire token_28_15;
    wire dep_chan_vld_29_15;
    wire [39:0] dep_chan_data_29_15;
    wire token_29_15;
    wire dep_chan_vld_30_15;
    wire [39:0] dep_chan_data_30_15;
    wire token_30_15;
    wire dep_chan_vld_31_15;
    wire [39:0] dep_chan_data_31_15;
    wire token_31_15;
    wire dep_chan_vld_32_15;
    wire [39:0] dep_chan_data_32_15;
    wire token_32_15;
    wire dep_chan_vld_33_15;
    wire [39:0] dep_chan_data_33_15;
    wire token_33_15;
    wire dep_chan_vld_34_15;
    wire [39:0] dep_chan_data_34_15;
    wire token_34_15;
    wire dep_chan_vld_35_15;
    wire [39:0] dep_chan_data_35_15;
    wire token_35_15;
    wire dep_chan_vld_36_15;
    wire [39:0] dep_chan_data_36_15;
    wire token_36_15;
    wire [32:0] proc_16_data_FIFO_blk;
    wire [32:0] proc_16_data_PIPO_blk;
    wire [32:0] proc_16_start_FIFO_blk;
    wire [32:0] proc_16_TLF_FIFO_blk;
    wire [32:0] proc_16_input_sync_blk;
    wire [32:0] proc_16_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_16;
    reg [32:0] proc_dep_vld_vec_16_reg;
    wire [32:0] in_chan_dep_vld_vec_16;
    wire [1319:0] in_chan_dep_data_vec_16;
    wire [32:0] token_in_vec_16;
    wire [32:0] out_chan_dep_vld_vec_16;
    wire [39:0] out_chan_dep_data_16;
    wire [32:0] token_out_vec_16;
    wire dl_detect_out_16;
    wire dep_chan_vld_0_16;
    wire [39:0] dep_chan_data_0_16;
    wire token_0_16;
    wire dep_chan_vld_1_16;
    wire [39:0] dep_chan_data_1_16;
    wire token_1_16;
    wire dep_chan_vld_3_16;
    wire [39:0] dep_chan_data_3_16;
    wire token_3_16;
    wire dep_chan_vld_6_16;
    wire [39:0] dep_chan_data_6_16;
    wire token_6_16;
    wire dep_chan_vld_7_16;
    wire [39:0] dep_chan_data_7_16;
    wire token_7_16;
    wire dep_chan_vld_8_16;
    wire [39:0] dep_chan_data_8_16;
    wire token_8_16;
    wire dep_chan_vld_9_16;
    wire [39:0] dep_chan_data_9_16;
    wire token_9_16;
    wire dep_chan_vld_10_16;
    wire [39:0] dep_chan_data_10_16;
    wire token_10_16;
    wire dep_chan_vld_11_16;
    wire [39:0] dep_chan_data_11_16;
    wire token_11_16;
    wire dep_chan_vld_12_16;
    wire [39:0] dep_chan_data_12_16;
    wire token_12_16;
    wire dep_chan_vld_13_16;
    wire [39:0] dep_chan_data_13_16;
    wire token_13_16;
    wire dep_chan_vld_14_16;
    wire [39:0] dep_chan_data_14_16;
    wire token_14_16;
    wire dep_chan_vld_15_16;
    wire [39:0] dep_chan_data_15_16;
    wire token_15_16;
    wire dep_chan_vld_17_16;
    wire [39:0] dep_chan_data_17_16;
    wire token_17_16;
    wire dep_chan_vld_18_16;
    wire [39:0] dep_chan_data_18_16;
    wire token_18_16;
    wire dep_chan_vld_19_16;
    wire [39:0] dep_chan_data_19_16;
    wire token_19_16;
    wire dep_chan_vld_20_16;
    wire [39:0] dep_chan_data_20_16;
    wire token_20_16;
    wire dep_chan_vld_21_16;
    wire [39:0] dep_chan_data_21_16;
    wire token_21_16;
    wire dep_chan_vld_22_16;
    wire [39:0] dep_chan_data_22_16;
    wire token_22_16;
    wire dep_chan_vld_23_16;
    wire [39:0] dep_chan_data_23_16;
    wire token_23_16;
    wire dep_chan_vld_24_16;
    wire [39:0] dep_chan_data_24_16;
    wire token_24_16;
    wire dep_chan_vld_25_16;
    wire [39:0] dep_chan_data_25_16;
    wire token_25_16;
    wire dep_chan_vld_26_16;
    wire [39:0] dep_chan_data_26_16;
    wire token_26_16;
    wire dep_chan_vld_27_16;
    wire [39:0] dep_chan_data_27_16;
    wire token_27_16;
    wire dep_chan_vld_28_16;
    wire [39:0] dep_chan_data_28_16;
    wire token_28_16;
    wire dep_chan_vld_29_16;
    wire [39:0] dep_chan_data_29_16;
    wire token_29_16;
    wire dep_chan_vld_30_16;
    wire [39:0] dep_chan_data_30_16;
    wire token_30_16;
    wire dep_chan_vld_31_16;
    wire [39:0] dep_chan_data_31_16;
    wire token_31_16;
    wire dep_chan_vld_32_16;
    wire [39:0] dep_chan_data_32_16;
    wire token_32_16;
    wire dep_chan_vld_33_16;
    wire [39:0] dep_chan_data_33_16;
    wire token_33_16;
    wire dep_chan_vld_34_16;
    wire [39:0] dep_chan_data_34_16;
    wire token_34_16;
    wire dep_chan_vld_35_16;
    wire [39:0] dep_chan_data_35_16;
    wire token_35_16;
    wire dep_chan_vld_36_16;
    wire [39:0] dep_chan_data_36_16;
    wire token_36_16;
    wire [32:0] proc_17_data_FIFO_blk;
    wire [32:0] proc_17_data_PIPO_blk;
    wire [32:0] proc_17_start_FIFO_blk;
    wire [32:0] proc_17_TLF_FIFO_blk;
    wire [32:0] proc_17_input_sync_blk;
    wire [32:0] proc_17_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_17;
    reg [32:0] proc_dep_vld_vec_17_reg;
    wire [32:0] in_chan_dep_vld_vec_17;
    wire [1319:0] in_chan_dep_data_vec_17;
    wire [32:0] token_in_vec_17;
    wire [32:0] out_chan_dep_vld_vec_17;
    wire [39:0] out_chan_dep_data_17;
    wire [32:0] token_out_vec_17;
    wire dl_detect_out_17;
    wire dep_chan_vld_0_17;
    wire [39:0] dep_chan_data_0_17;
    wire token_0_17;
    wire dep_chan_vld_1_17;
    wire [39:0] dep_chan_data_1_17;
    wire token_1_17;
    wire dep_chan_vld_3_17;
    wire [39:0] dep_chan_data_3_17;
    wire token_3_17;
    wire dep_chan_vld_6_17;
    wire [39:0] dep_chan_data_6_17;
    wire token_6_17;
    wire dep_chan_vld_7_17;
    wire [39:0] dep_chan_data_7_17;
    wire token_7_17;
    wire dep_chan_vld_8_17;
    wire [39:0] dep_chan_data_8_17;
    wire token_8_17;
    wire dep_chan_vld_9_17;
    wire [39:0] dep_chan_data_9_17;
    wire token_9_17;
    wire dep_chan_vld_10_17;
    wire [39:0] dep_chan_data_10_17;
    wire token_10_17;
    wire dep_chan_vld_11_17;
    wire [39:0] dep_chan_data_11_17;
    wire token_11_17;
    wire dep_chan_vld_12_17;
    wire [39:0] dep_chan_data_12_17;
    wire token_12_17;
    wire dep_chan_vld_13_17;
    wire [39:0] dep_chan_data_13_17;
    wire token_13_17;
    wire dep_chan_vld_14_17;
    wire [39:0] dep_chan_data_14_17;
    wire token_14_17;
    wire dep_chan_vld_15_17;
    wire [39:0] dep_chan_data_15_17;
    wire token_15_17;
    wire dep_chan_vld_16_17;
    wire [39:0] dep_chan_data_16_17;
    wire token_16_17;
    wire dep_chan_vld_18_17;
    wire [39:0] dep_chan_data_18_17;
    wire token_18_17;
    wire dep_chan_vld_19_17;
    wire [39:0] dep_chan_data_19_17;
    wire token_19_17;
    wire dep_chan_vld_20_17;
    wire [39:0] dep_chan_data_20_17;
    wire token_20_17;
    wire dep_chan_vld_21_17;
    wire [39:0] dep_chan_data_21_17;
    wire token_21_17;
    wire dep_chan_vld_22_17;
    wire [39:0] dep_chan_data_22_17;
    wire token_22_17;
    wire dep_chan_vld_23_17;
    wire [39:0] dep_chan_data_23_17;
    wire token_23_17;
    wire dep_chan_vld_24_17;
    wire [39:0] dep_chan_data_24_17;
    wire token_24_17;
    wire dep_chan_vld_25_17;
    wire [39:0] dep_chan_data_25_17;
    wire token_25_17;
    wire dep_chan_vld_26_17;
    wire [39:0] dep_chan_data_26_17;
    wire token_26_17;
    wire dep_chan_vld_27_17;
    wire [39:0] dep_chan_data_27_17;
    wire token_27_17;
    wire dep_chan_vld_28_17;
    wire [39:0] dep_chan_data_28_17;
    wire token_28_17;
    wire dep_chan_vld_29_17;
    wire [39:0] dep_chan_data_29_17;
    wire token_29_17;
    wire dep_chan_vld_30_17;
    wire [39:0] dep_chan_data_30_17;
    wire token_30_17;
    wire dep_chan_vld_31_17;
    wire [39:0] dep_chan_data_31_17;
    wire token_31_17;
    wire dep_chan_vld_32_17;
    wire [39:0] dep_chan_data_32_17;
    wire token_32_17;
    wire dep_chan_vld_33_17;
    wire [39:0] dep_chan_data_33_17;
    wire token_33_17;
    wire dep_chan_vld_34_17;
    wire [39:0] dep_chan_data_34_17;
    wire token_34_17;
    wire dep_chan_vld_35_17;
    wire [39:0] dep_chan_data_35_17;
    wire token_35_17;
    wire dep_chan_vld_36_17;
    wire [39:0] dep_chan_data_36_17;
    wire token_36_17;
    wire [32:0] proc_18_data_FIFO_blk;
    wire [32:0] proc_18_data_PIPO_blk;
    wire [32:0] proc_18_start_FIFO_blk;
    wire [32:0] proc_18_TLF_FIFO_blk;
    wire [32:0] proc_18_input_sync_blk;
    wire [32:0] proc_18_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_18;
    reg [32:0] proc_dep_vld_vec_18_reg;
    wire [32:0] in_chan_dep_vld_vec_18;
    wire [1319:0] in_chan_dep_data_vec_18;
    wire [32:0] token_in_vec_18;
    wire [32:0] out_chan_dep_vld_vec_18;
    wire [39:0] out_chan_dep_data_18;
    wire [32:0] token_out_vec_18;
    wire dl_detect_out_18;
    wire dep_chan_vld_0_18;
    wire [39:0] dep_chan_data_0_18;
    wire token_0_18;
    wire dep_chan_vld_1_18;
    wire [39:0] dep_chan_data_1_18;
    wire token_1_18;
    wire dep_chan_vld_3_18;
    wire [39:0] dep_chan_data_3_18;
    wire token_3_18;
    wire dep_chan_vld_6_18;
    wire [39:0] dep_chan_data_6_18;
    wire token_6_18;
    wire dep_chan_vld_7_18;
    wire [39:0] dep_chan_data_7_18;
    wire token_7_18;
    wire dep_chan_vld_8_18;
    wire [39:0] dep_chan_data_8_18;
    wire token_8_18;
    wire dep_chan_vld_9_18;
    wire [39:0] dep_chan_data_9_18;
    wire token_9_18;
    wire dep_chan_vld_10_18;
    wire [39:0] dep_chan_data_10_18;
    wire token_10_18;
    wire dep_chan_vld_11_18;
    wire [39:0] dep_chan_data_11_18;
    wire token_11_18;
    wire dep_chan_vld_12_18;
    wire [39:0] dep_chan_data_12_18;
    wire token_12_18;
    wire dep_chan_vld_13_18;
    wire [39:0] dep_chan_data_13_18;
    wire token_13_18;
    wire dep_chan_vld_14_18;
    wire [39:0] dep_chan_data_14_18;
    wire token_14_18;
    wire dep_chan_vld_15_18;
    wire [39:0] dep_chan_data_15_18;
    wire token_15_18;
    wire dep_chan_vld_16_18;
    wire [39:0] dep_chan_data_16_18;
    wire token_16_18;
    wire dep_chan_vld_17_18;
    wire [39:0] dep_chan_data_17_18;
    wire token_17_18;
    wire dep_chan_vld_19_18;
    wire [39:0] dep_chan_data_19_18;
    wire token_19_18;
    wire dep_chan_vld_20_18;
    wire [39:0] dep_chan_data_20_18;
    wire token_20_18;
    wire dep_chan_vld_21_18;
    wire [39:0] dep_chan_data_21_18;
    wire token_21_18;
    wire dep_chan_vld_22_18;
    wire [39:0] dep_chan_data_22_18;
    wire token_22_18;
    wire dep_chan_vld_23_18;
    wire [39:0] dep_chan_data_23_18;
    wire token_23_18;
    wire dep_chan_vld_24_18;
    wire [39:0] dep_chan_data_24_18;
    wire token_24_18;
    wire dep_chan_vld_25_18;
    wire [39:0] dep_chan_data_25_18;
    wire token_25_18;
    wire dep_chan_vld_26_18;
    wire [39:0] dep_chan_data_26_18;
    wire token_26_18;
    wire dep_chan_vld_27_18;
    wire [39:0] dep_chan_data_27_18;
    wire token_27_18;
    wire dep_chan_vld_28_18;
    wire [39:0] dep_chan_data_28_18;
    wire token_28_18;
    wire dep_chan_vld_29_18;
    wire [39:0] dep_chan_data_29_18;
    wire token_29_18;
    wire dep_chan_vld_30_18;
    wire [39:0] dep_chan_data_30_18;
    wire token_30_18;
    wire dep_chan_vld_31_18;
    wire [39:0] dep_chan_data_31_18;
    wire token_31_18;
    wire dep_chan_vld_32_18;
    wire [39:0] dep_chan_data_32_18;
    wire token_32_18;
    wire dep_chan_vld_33_18;
    wire [39:0] dep_chan_data_33_18;
    wire token_33_18;
    wire dep_chan_vld_34_18;
    wire [39:0] dep_chan_data_34_18;
    wire token_34_18;
    wire dep_chan_vld_35_18;
    wire [39:0] dep_chan_data_35_18;
    wire token_35_18;
    wire dep_chan_vld_36_18;
    wire [39:0] dep_chan_data_36_18;
    wire token_36_18;
    wire [32:0] proc_19_data_FIFO_blk;
    wire [32:0] proc_19_data_PIPO_blk;
    wire [32:0] proc_19_start_FIFO_blk;
    wire [32:0] proc_19_TLF_FIFO_blk;
    wire [32:0] proc_19_input_sync_blk;
    wire [32:0] proc_19_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_19;
    reg [32:0] proc_dep_vld_vec_19_reg;
    wire [32:0] in_chan_dep_vld_vec_19;
    wire [1319:0] in_chan_dep_data_vec_19;
    wire [32:0] token_in_vec_19;
    wire [32:0] out_chan_dep_vld_vec_19;
    wire [39:0] out_chan_dep_data_19;
    wire [32:0] token_out_vec_19;
    wire dl_detect_out_19;
    wire dep_chan_vld_0_19;
    wire [39:0] dep_chan_data_0_19;
    wire token_0_19;
    wire dep_chan_vld_1_19;
    wire [39:0] dep_chan_data_1_19;
    wire token_1_19;
    wire dep_chan_vld_3_19;
    wire [39:0] dep_chan_data_3_19;
    wire token_3_19;
    wire dep_chan_vld_6_19;
    wire [39:0] dep_chan_data_6_19;
    wire token_6_19;
    wire dep_chan_vld_7_19;
    wire [39:0] dep_chan_data_7_19;
    wire token_7_19;
    wire dep_chan_vld_8_19;
    wire [39:0] dep_chan_data_8_19;
    wire token_8_19;
    wire dep_chan_vld_9_19;
    wire [39:0] dep_chan_data_9_19;
    wire token_9_19;
    wire dep_chan_vld_10_19;
    wire [39:0] dep_chan_data_10_19;
    wire token_10_19;
    wire dep_chan_vld_11_19;
    wire [39:0] dep_chan_data_11_19;
    wire token_11_19;
    wire dep_chan_vld_12_19;
    wire [39:0] dep_chan_data_12_19;
    wire token_12_19;
    wire dep_chan_vld_13_19;
    wire [39:0] dep_chan_data_13_19;
    wire token_13_19;
    wire dep_chan_vld_14_19;
    wire [39:0] dep_chan_data_14_19;
    wire token_14_19;
    wire dep_chan_vld_15_19;
    wire [39:0] dep_chan_data_15_19;
    wire token_15_19;
    wire dep_chan_vld_16_19;
    wire [39:0] dep_chan_data_16_19;
    wire token_16_19;
    wire dep_chan_vld_17_19;
    wire [39:0] dep_chan_data_17_19;
    wire token_17_19;
    wire dep_chan_vld_18_19;
    wire [39:0] dep_chan_data_18_19;
    wire token_18_19;
    wire dep_chan_vld_20_19;
    wire [39:0] dep_chan_data_20_19;
    wire token_20_19;
    wire dep_chan_vld_21_19;
    wire [39:0] dep_chan_data_21_19;
    wire token_21_19;
    wire dep_chan_vld_22_19;
    wire [39:0] dep_chan_data_22_19;
    wire token_22_19;
    wire dep_chan_vld_23_19;
    wire [39:0] dep_chan_data_23_19;
    wire token_23_19;
    wire dep_chan_vld_24_19;
    wire [39:0] dep_chan_data_24_19;
    wire token_24_19;
    wire dep_chan_vld_25_19;
    wire [39:0] dep_chan_data_25_19;
    wire token_25_19;
    wire dep_chan_vld_26_19;
    wire [39:0] dep_chan_data_26_19;
    wire token_26_19;
    wire dep_chan_vld_27_19;
    wire [39:0] dep_chan_data_27_19;
    wire token_27_19;
    wire dep_chan_vld_28_19;
    wire [39:0] dep_chan_data_28_19;
    wire token_28_19;
    wire dep_chan_vld_29_19;
    wire [39:0] dep_chan_data_29_19;
    wire token_29_19;
    wire dep_chan_vld_30_19;
    wire [39:0] dep_chan_data_30_19;
    wire token_30_19;
    wire dep_chan_vld_31_19;
    wire [39:0] dep_chan_data_31_19;
    wire token_31_19;
    wire dep_chan_vld_32_19;
    wire [39:0] dep_chan_data_32_19;
    wire token_32_19;
    wire dep_chan_vld_33_19;
    wire [39:0] dep_chan_data_33_19;
    wire token_33_19;
    wire dep_chan_vld_34_19;
    wire [39:0] dep_chan_data_34_19;
    wire token_34_19;
    wire dep_chan_vld_35_19;
    wire [39:0] dep_chan_data_35_19;
    wire token_35_19;
    wire dep_chan_vld_36_19;
    wire [39:0] dep_chan_data_36_19;
    wire token_36_19;
    wire [32:0] proc_20_data_FIFO_blk;
    wire [32:0] proc_20_data_PIPO_blk;
    wire [32:0] proc_20_start_FIFO_blk;
    wire [32:0] proc_20_TLF_FIFO_blk;
    wire [32:0] proc_20_input_sync_blk;
    wire [32:0] proc_20_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_20;
    reg [32:0] proc_dep_vld_vec_20_reg;
    wire [32:0] in_chan_dep_vld_vec_20;
    wire [1319:0] in_chan_dep_data_vec_20;
    wire [32:0] token_in_vec_20;
    wire [32:0] out_chan_dep_vld_vec_20;
    wire [39:0] out_chan_dep_data_20;
    wire [32:0] token_out_vec_20;
    wire dl_detect_out_20;
    wire dep_chan_vld_0_20;
    wire [39:0] dep_chan_data_0_20;
    wire token_0_20;
    wire dep_chan_vld_1_20;
    wire [39:0] dep_chan_data_1_20;
    wire token_1_20;
    wire dep_chan_vld_3_20;
    wire [39:0] dep_chan_data_3_20;
    wire token_3_20;
    wire dep_chan_vld_6_20;
    wire [39:0] dep_chan_data_6_20;
    wire token_6_20;
    wire dep_chan_vld_7_20;
    wire [39:0] dep_chan_data_7_20;
    wire token_7_20;
    wire dep_chan_vld_8_20;
    wire [39:0] dep_chan_data_8_20;
    wire token_8_20;
    wire dep_chan_vld_9_20;
    wire [39:0] dep_chan_data_9_20;
    wire token_9_20;
    wire dep_chan_vld_10_20;
    wire [39:0] dep_chan_data_10_20;
    wire token_10_20;
    wire dep_chan_vld_11_20;
    wire [39:0] dep_chan_data_11_20;
    wire token_11_20;
    wire dep_chan_vld_12_20;
    wire [39:0] dep_chan_data_12_20;
    wire token_12_20;
    wire dep_chan_vld_13_20;
    wire [39:0] dep_chan_data_13_20;
    wire token_13_20;
    wire dep_chan_vld_14_20;
    wire [39:0] dep_chan_data_14_20;
    wire token_14_20;
    wire dep_chan_vld_15_20;
    wire [39:0] dep_chan_data_15_20;
    wire token_15_20;
    wire dep_chan_vld_16_20;
    wire [39:0] dep_chan_data_16_20;
    wire token_16_20;
    wire dep_chan_vld_17_20;
    wire [39:0] dep_chan_data_17_20;
    wire token_17_20;
    wire dep_chan_vld_18_20;
    wire [39:0] dep_chan_data_18_20;
    wire token_18_20;
    wire dep_chan_vld_19_20;
    wire [39:0] dep_chan_data_19_20;
    wire token_19_20;
    wire dep_chan_vld_21_20;
    wire [39:0] dep_chan_data_21_20;
    wire token_21_20;
    wire dep_chan_vld_22_20;
    wire [39:0] dep_chan_data_22_20;
    wire token_22_20;
    wire dep_chan_vld_23_20;
    wire [39:0] dep_chan_data_23_20;
    wire token_23_20;
    wire dep_chan_vld_24_20;
    wire [39:0] dep_chan_data_24_20;
    wire token_24_20;
    wire dep_chan_vld_25_20;
    wire [39:0] dep_chan_data_25_20;
    wire token_25_20;
    wire dep_chan_vld_26_20;
    wire [39:0] dep_chan_data_26_20;
    wire token_26_20;
    wire dep_chan_vld_27_20;
    wire [39:0] dep_chan_data_27_20;
    wire token_27_20;
    wire dep_chan_vld_28_20;
    wire [39:0] dep_chan_data_28_20;
    wire token_28_20;
    wire dep_chan_vld_29_20;
    wire [39:0] dep_chan_data_29_20;
    wire token_29_20;
    wire dep_chan_vld_30_20;
    wire [39:0] dep_chan_data_30_20;
    wire token_30_20;
    wire dep_chan_vld_31_20;
    wire [39:0] dep_chan_data_31_20;
    wire token_31_20;
    wire dep_chan_vld_32_20;
    wire [39:0] dep_chan_data_32_20;
    wire token_32_20;
    wire dep_chan_vld_33_20;
    wire [39:0] dep_chan_data_33_20;
    wire token_33_20;
    wire dep_chan_vld_34_20;
    wire [39:0] dep_chan_data_34_20;
    wire token_34_20;
    wire dep_chan_vld_35_20;
    wire [39:0] dep_chan_data_35_20;
    wire token_35_20;
    wire dep_chan_vld_36_20;
    wire [39:0] dep_chan_data_36_20;
    wire token_36_20;
    wire [32:0] proc_21_data_FIFO_blk;
    wire [32:0] proc_21_data_PIPO_blk;
    wire [32:0] proc_21_start_FIFO_blk;
    wire [32:0] proc_21_TLF_FIFO_blk;
    wire [32:0] proc_21_input_sync_blk;
    wire [32:0] proc_21_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_21;
    reg [32:0] proc_dep_vld_vec_21_reg;
    wire [32:0] in_chan_dep_vld_vec_21;
    wire [1319:0] in_chan_dep_data_vec_21;
    wire [32:0] token_in_vec_21;
    wire [32:0] out_chan_dep_vld_vec_21;
    wire [39:0] out_chan_dep_data_21;
    wire [32:0] token_out_vec_21;
    wire dl_detect_out_21;
    wire dep_chan_vld_0_21;
    wire [39:0] dep_chan_data_0_21;
    wire token_0_21;
    wire dep_chan_vld_1_21;
    wire [39:0] dep_chan_data_1_21;
    wire token_1_21;
    wire dep_chan_vld_3_21;
    wire [39:0] dep_chan_data_3_21;
    wire token_3_21;
    wire dep_chan_vld_6_21;
    wire [39:0] dep_chan_data_6_21;
    wire token_6_21;
    wire dep_chan_vld_7_21;
    wire [39:0] dep_chan_data_7_21;
    wire token_7_21;
    wire dep_chan_vld_8_21;
    wire [39:0] dep_chan_data_8_21;
    wire token_8_21;
    wire dep_chan_vld_9_21;
    wire [39:0] dep_chan_data_9_21;
    wire token_9_21;
    wire dep_chan_vld_10_21;
    wire [39:0] dep_chan_data_10_21;
    wire token_10_21;
    wire dep_chan_vld_11_21;
    wire [39:0] dep_chan_data_11_21;
    wire token_11_21;
    wire dep_chan_vld_12_21;
    wire [39:0] dep_chan_data_12_21;
    wire token_12_21;
    wire dep_chan_vld_13_21;
    wire [39:0] dep_chan_data_13_21;
    wire token_13_21;
    wire dep_chan_vld_14_21;
    wire [39:0] dep_chan_data_14_21;
    wire token_14_21;
    wire dep_chan_vld_15_21;
    wire [39:0] dep_chan_data_15_21;
    wire token_15_21;
    wire dep_chan_vld_16_21;
    wire [39:0] dep_chan_data_16_21;
    wire token_16_21;
    wire dep_chan_vld_17_21;
    wire [39:0] dep_chan_data_17_21;
    wire token_17_21;
    wire dep_chan_vld_18_21;
    wire [39:0] dep_chan_data_18_21;
    wire token_18_21;
    wire dep_chan_vld_19_21;
    wire [39:0] dep_chan_data_19_21;
    wire token_19_21;
    wire dep_chan_vld_20_21;
    wire [39:0] dep_chan_data_20_21;
    wire token_20_21;
    wire dep_chan_vld_22_21;
    wire [39:0] dep_chan_data_22_21;
    wire token_22_21;
    wire dep_chan_vld_23_21;
    wire [39:0] dep_chan_data_23_21;
    wire token_23_21;
    wire dep_chan_vld_24_21;
    wire [39:0] dep_chan_data_24_21;
    wire token_24_21;
    wire dep_chan_vld_25_21;
    wire [39:0] dep_chan_data_25_21;
    wire token_25_21;
    wire dep_chan_vld_26_21;
    wire [39:0] dep_chan_data_26_21;
    wire token_26_21;
    wire dep_chan_vld_27_21;
    wire [39:0] dep_chan_data_27_21;
    wire token_27_21;
    wire dep_chan_vld_28_21;
    wire [39:0] dep_chan_data_28_21;
    wire token_28_21;
    wire dep_chan_vld_29_21;
    wire [39:0] dep_chan_data_29_21;
    wire token_29_21;
    wire dep_chan_vld_30_21;
    wire [39:0] dep_chan_data_30_21;
    wire token_30_21;
    wire dep_chan_vld_31_21;
    wire [39:0] dep_chan_data_31_21;
    wire token_31_21;
    wire dep_chan_vld_32_21;
    wire [39:0] dep_chan_data_32_21;
    wire token_32_21;
    wire dep_chan_vld_33_21;
    wire [39:0] dep_chan_data_33_21;
    wire token_33_21;
    wire dep_chan_vld_34_21;
    wire [39:0] dep_chan_data_34_21;
    wire token_34_21;
    wire dep_chan_vld_35_21;
    wire [39:0] dep_chan_data_35_21;
    wire token_35_21;
    wire dep_chan_vld_36_21;
    wire [39:0] dep_chan_data_36_21;
    wire token_36_21;
    wire [32:0] proc_22_data_FIFO_blk;
    wire [32:0] proc_22_data_PIPO_blk;
    wire [32:0] proc_22_start_FIFO_blk;
    wire [32:0] proc_22_TLF_FIFO_blk;
    wire [32:0] proc_22_input_sync_blk;
    wire [32:0] proc_22_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_22;
    reg [32:0] proc_dep_vld_vec_22_reg;
    wire [32:0] in_chan_dep_vld_vec_22;
    wire [1319:0] in_chan_dep_data_vec_22;
    wire [32:0] token_in_vec_22;
    wire [32:0] out_chan_dep_vld_vec_22;
    wire [39:0] out_chan_dep_data_22;
    wire [32:0] token_out_vec_22;
    wire dl_detect_out_22;
    wire dep_chan_vld_0_22;
    wire [39:0] dep_chan_data_0_22;
    wire token_0_22;
    wire dep_chan_vld_1_22;
    wire [39:0] dep_chan_data_1_22;
    wire token_1_22;
    wire dep_chan_vld_3_22;
    wire [39:0] dep_chan_data_3_22;
    wire token_3_22;
    wire dep_chan_vld_6_22;
    wire [39:0] dep_chan_data_6_22;
    wire token_6_22;
    wire dep_chan_vld_7_22;
    wire [39:0] dep_chan_data_7_22;
    wire token_7_22;
    wire dep_chan_vld_8_22;
    wire [39:0] dep_chan_data_8_22;
    wire token_8_22;
    wire dep_chan_vld_9_22;
    wire [39:0] dep_chan_data_9_22;
    wire token_9_22;
    wire dep_chan_vld_10_22;
    wire [39:0] dep_chan_data_10_22;
    wire token_10_22;
    wire dep_chan_vld_11_22;
    wire [39:0] dep_chan_data_11_22;
    wire token_11_22;
    wire dep_chan_vld_12_22;
    wire [39:0] dep_chan_data_12_22;
    wire token_12_22;
    wire dep_chan_vld_13_22;
    wire [39:0] dep_chan_data_13_22;
    wire token_13_22;
    wire dep_chan_vld_14_22;
    wire [39:0] dep_chan_data_14_22;
    wire token_14_22;
    wire dep_chan_vld_15_22;
    wire [39:0] dep_chan_data_15_22;
    wire token_15_22;
    wire dep_chan_vld_16_22;
    wire [39:0] dep_chan_data_16_22;
    wire token_16_22;
    wire dep_chan_vld_17_22;
    wire [39:0] dep_chan_data_17_22;
    wire token_17_22;
    wire dep_chan_vld_18_22;
    wire [39:0] dep_chan_data_18_22;
    wire token_18_22;
    wire dep_chan_vld_19_22;
    wire [39:0] dep_chan_data_19_22;
    wire token_19_22;
    wire dep_chan_vld_20_22;
    wire [39:0] dep_chan_data_20_22;
    wire token_20_22;
    wire dep_chan_vld_21_22;
    wire [39:0] dep_chan_data_21_22;
    wire token_21_22;
    wire dep_chan_vld_23_22;
    wire [39:0] dep_chan_data_23_22;
    wire token_23_22;
    wire dep_chan_vld_24_22;
    wire [39:0] dep_chan_data_24_22;
    wire token_24_22;
    wire dep_chan_vld_25_22;
    wire [39:0] dep_chan_data_25_22;
    wire token_25_22;
    wire dep_chan_vld_26_22;
    wire [39:0] dep_chan_data_26_22;
    wire token_26_22;
    wire dep_chan_vld_27_22;
    wire [39:0] dep_chan_data_27_22;
    wire token_27_22;
    wire dep_chan_vld_28_22;
    wire [39:0] dep_chan_data_28_22;
    wire token_28_22;
    wire dep_chan_vld_29_22;
    wire [39:0] dep_chan_data_29_22;
    wire token_29_22;
    wire dep_chan_vld_30_22;
    wire [39:0] dep_chan_data_30_22;
    wire token_30_22;
    wire dep_chan_vld_31_22;
    wire [39:0] dep_chan_data_31_22;
    wire token_31_22;
    wire dep_chan_vld_32_22;
    wire [39:0] dep_chan_data_32_22;
    wire token_32_22;
    wire dep_chan_vld_33_22;
    wire [39:0] dep_chan_data_33_22;
    wire token_33_22;
    wire dep_chan_vld_34_22;
    wire [39:0] dep_chan_data_34_22;
    wire token_34_22;
    wire dep_chan_vld_35_22;
    wire [39:0] dep_chan_data_35_22;
    wire token_35_22;
    wire dep_chan_vld_36_22;
    wire [39:0] dep_chan_data_36_22;
    wire token_36_22;
    wire [32:0] proc_23_data_FIFO_blk;
    wire [32:0] proc_23_data_PIPO_blk;
    wire [32:0] proc_23_start_FIFO_blk;
    wire [32:0] proc_23_TLF_FIFO_blk;
    wire [32:0] proc_23_input_sync_blk;
    wire [32:0] proc_23_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_23;
    reg [32:0] proc_dep_vld_vec_23_reg;
    wire [32:0] in_chan_dep_vld_vec_23;
    wire [1319:0] in_chan_dep_data_vec_23;
    wire [32:0] token_in_vec_23;
    wire [32:0] out_chan_dep_vld_vec_23;
    wire [39:0] out_chan_dep_data_23;
    wire [32:0] token_out_vec_23;
    wire dl_detect_out_23;
    wire dep_chan_vld_0_23;
    wire [39:0] dep_chan_data_0_23;
    wire token_0_23;
    wire dep_chan_vld_1_23;
    wire [39:0] dep_chan_data_1_23;
    wire token_1_23;
    wire dep_chan_vld_3_23;
    wire [39:0] dep_chan_data_3_23;
    wire token_3_23;
    wire dep_chan_vld_6_23;
    wire [39:0] dep_chan_data_6_23;
    wire token_6_23;
    wire dep_chan_vld_7_23;
    wire [39:0] dep_chan_data_7_23;
    wire token_7_23;
    wire dep_chan_vld_8_23;
    wire [39:0] dep_chan_data_8_23;
    wire token_8_23;
    wire dep_chan_vld_9_23;
    wire [39:0] dep_chan_data_9_23;
    wire token_9_23;
    wire dep_chan_vld_10_23;
    wire [39:0] dep_chan_data_10_23;
    wire token_10_23;
    wire dep_chan_vld_11_23;
    wire [39:0] dep_chan_data_11_23;
    wire token_11_23;
    wire dep_chan_vld_12_23;
    wire [39:0] dep_chan_data_12_23;
    wire token_12_23;
    wire dep_chan_vld_13_23;
    wire [39:0] dep_chan_data_13_23;
    wire token_13_23;
    wire dep_chan_vld_14_23;
    wire [39:0] dep_chan_data_14_23;
    wire token_14_23;
    wire dep_chan_vld_15_23;
    wire [39:0] dep_chan_data_15_23;
    wire token_15_23;
    wire dep_chan_vld_16_23;
    wire [39:0] dep_chan_data_16_23;
    wire token_16_23;
    wire dep_chan_vld_17_23;
    wire [39:0] dep_chan_data_17_23;
    wire token_17_23;
    wire dep_chan_vld_18_23;
    wire [39:0] dep_chan_data_18_23;
    wire token_18_23;
    wire dep_chan_vld_19_23;
    wire [39:0] dep_chan_data_19_23;
    wire token_19_23;
    wire dep_chan_vld_20_23;
    wire [39:0] dep_chan_data_20_23;
    wire token_20_23;
    wire dep_chan_vld_21_23;
    wire [39:0] dep_chan_data_21_23;
    wire token_21_23;
    wire dep_chan_vld_22_23;
    wire [39:0] dep_chan_data_22_23;
    wire token_22_23;
    wire dep_chan_vld_24_23;
    wire [39:0] dep_chan_data_24_23;
    wire token_24_23;
    wire dep_chan_vld_25_23;
    wire [39:0] dep_chan_data_25_23;
    wire token_25_23;
    wire dep_chan_vld_26_23;
    wire [39:0] dep_chan_data_26_23;
    wire token_26_23;
    wire dep_chan_vld_27_23;
    wire [39:0] dep_chan_data_27_23;
    wire token_27_23;
    wire dep_chan_vld_28_23;
    wire [39:0] dep_chan_data_28_23;
    wire token_28_23;
    wire dep_chan_vld_29_23;
    wire [39:0] dep_chan_data_29_23;
    wire token_29_23;
    wire dep_chan_vld_30_23;
    wire [39:0] dep_chan_data_30_23;
    wire token_30_23;
    wire dep_chan_vld_31_23;
    wire [39:0] dep_chan_data_31_23;
    wire token_31_23;
    wire dep_chan_vld_32_23;
    wire [39:0] dep_chan_data_32_23;
    wire token_32_23;
    wire dep_chan_vld_33_23;
    wire [39:0] dep_chan_data_33_23;
    wire token_33_23;
    wire dep_chan_vld_34_23;
    wire [39:0] dep_chan_data_34_23;
    wire token_34_23;
    wire dep_chan_vld_35_23;
    wire [39:0] dep_chan_data_35_23;
    wire token_35_23;
    wire dep_chan_vld_36_23;
    wire [39:0] dep_chan_data_36_23;
    wire token_36_23;
    wire [32:0] proc_24_data_FIFO_blk;
    wire [32:0] proc_24_data_PIPO_blk;
    wire [32:0] proc_24_start_FIFO_blk;
    wire [32:0] proc_24_TLF_FIFO_blk;
    wire [32:0] proc_24_input_sync_blk;
    wire [32:0] proc_24_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_24;
    reg [32:0] proc_dep_vld_vec_24_reg;
    wire [32:0] in_chan_dep_vld_vec_24;
    wire [1319:0] in_chan_dep_data_vec_24;
    wire [32:0] token_in_vec_24;
    wire [32:0] out_chan_dep_vld_vec_24;
    wire [39:0] out_chan_dep_data_24;
    wire [32:0] token_out_vec_24;
    wire dl_detect_out_24;
    wire dep_chan_vld_0_24;
    wire [39:0] dep_chan_data_0_24;
    wire token_0_24;
    wire dep_chan_vld_1_24;
    wire [39:0] dep_chan_data_1_24;
    wire token_1_24;
    wire dep_chan_vld_3_24;
    wire [39:0] dep_chan_data_3_24;
    wire token_3_24;
    wire dep_chan_vld_6_24;
    wire [39:0] dep_chan_data_6_24;
    wire token_6_24;
    wire dep_chan_vld_7_24;
    wire [39:0] dep_chan_data_7_24;
    wire token_7_24;
    wire dep_chan_vld_8_24;
    wire [39:0] dep_chan_data_8_24;
    wire token_8_24;
    wire dep_chan_vld_9_24;
    wire [39:0] dep_chan_data_9_24;
    wire token_9_24;
    wire dep_chan_vld_10_24;
    wire [39:0] dep_chan_data_10_24;
    wire token_10_24;
    wire dep_chan_vld_11_24;
    wire [39:0] dep_chan_data_11_24;
    wire token_11_24;
    wire dep_chan_vld_12_24;
    wire [39:0] dep_chan_data_12_24;
    wire token_12_24;
    wire dep_chan_vld_13_24;
    wire [39:0] dep_chan_data_13_24;
    wire token_13_24;
    wire dep_chan_vld_14_24;
    wire [39:0] dep_chan_data_14_24;
    wire token_14_24;
    wire dep_chan_vld_15_24;
    wire [39:0] dep_chan_data_15_24;
    wire token_15_24;
    wire dep_chan_vld_16_24;
    wire [39:0] dep_chan_data_16_24;
    wire token_16_24;
    wire dep_chan_vld_17_24;
    wire [39:0] dep_chan_data_17_24;
    wire token_17_24;
    wire dep_chan_vld_18_24;
    wire [39:0] dep_chan_data_18_24;
    wire token_18_24;
    wire dep_chan_vld_19_24;
    wire [39:0] dep_chan_data_19_24;
    wire token_19_24;
    wire dep_chan_vld_20_24;
    wire [39:0] dep_chan_data_20_24;
    wire token_20_24;
    wire dep_chan_vld_21_24;
    wire [39:0] dep_chan_data_21_24;
    wire token_21_24;
    wire dep_chan_vld_22_24;
    wire [39:0] dep_chan_data_22_24;
    wire token_22_24;
    wire dep_chan_vld_23_24;
    wire [39:0] dep_chan_data_23_24;
    wire token_23_24;
    wire dep_chan_vld_25_24;
    wire [39:0] dep_chan_data_25_24;
    wire token_25_24;
    wire dep_chan_vld_26_24;
    wire [39:0] dep_chan_data_26_24;
    wire token_26_24;
    wire dep_chan_vld_27_24;
    wire [39:0] dep_chan_data_27_24;
    wire token_27_24;
    wire dep_chan_vld_28_24;
    wire [39:0] dep_chan_data_28_24;
    wire token_28_24;
    wire dep_chan_vld_29_24;
    wire [39:0] dep_chan_data_29_24;
    wire token_29_24;
    wire dep_chan_vld_30_24;
    wire [39:0] dep_chan_data_30_24;
    wire token_30_24;
    wire dep_chan_vld_31_24;
    wire [39:0] dep_chan_data_31_24;
    wire token_31_24;
    wire dep_chan_vld_32_24;
    wire [39:0] dep_chan_data_32_24;
    wire token_32_24;
    wire dep_chan_vld_33_24;
    wire [39:0] dep_chan_data_33_24;
    wire token_33_24;
    wire dep_chan_vld_34_24;
    wire [39:0] dep_chan_data_34_24;
    wire token_34_24;
    wire dep_chan_vld_35_24;
    wire [39:0] dep_chan_data_35_24;
    wire token_35_24;
    wire dep_chan_vld_36_24;
    wire [39:0] dep_chan_data_36_24;
    wire token_36_24;
    wire [32:0] proc_25_data_FIFO_blk;
    wire [32:0] proc_25_data_PIPO_blk;
    wire [32:0] proc_25_start_FIFO_blk;
    wire [32:0] proc_25_TLF_FIFO_blk;
    wire [32:0] proc_25_input_sync_blk;
    wire [32:0] proc_25_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_25;
    reg [32:0] proc_dep_vld_vec_25_reg;
    wire [32:0] in_chan_dep_vld_vec_25;
    wire [1319:0] in_chan_dep_data_vec_25;
    wire [32:0] token_in_vec_25;
    wire [32:0] out_chan_dep_vld_vec_25;
    wire [39:0] out_chan_dep_data_25;
    wire [32:0] token_out_vec_25;
    wire dl_detect_out_25;
    wire dep_chan_vld_0_25;
    wire [39:0] dep_chan_data_0_25;
    wire token_0_25;
    wire dep_chan_vld_1_25;
    wire [39:0] dep_chan_data_1_25;
    wire token_1_25;
    wire dep_chan_vld_3_25;
    wire [39:0] dep_chan_data_3_25;
    wire token_3_25;
    wire dep_chan_vld_6_25;
    wire [39:0] dep_chan_data_6_25;
    wire token_6_25;
    wire dep_chan_vld_7_25;
    wire [39:0] dep_chan_data_7_25;
    wire token_7_25;
    wire dep_chan_vld_8_25;
    wire [39:0] dep_chan_data_8_25;
    wire token_8_25;
    wire dep_chan_vld_9_25;
    wire [39:0] dep_chan_data_9_25;
    wire token_9_25;
    wire dep_chan_vld_10_25;
    wire [39:0] dep_chan_data_10_25;
    wire token_10_25;
    wire dep_chan_vld_11_25;
    wire [39:0] dep_chan_data_11_25;
    wire token_11_25;
    wire dep_chan_vld_12_25;
    wire [39:0] dep_chan_data_12_25;
    wire token_12_25;
    wire dep_chan_vld_13_25;
    wire [39:0] dep_chan_data_13_25;
    wire token_13_25;
    wire dep_chan_vld_14_25;
    wire [39:0] dep_chan_data_14_25;
    wire token_14_25;
    wire dep_chan_vld_15_25;
    wire [39:0] dep_chan_data_15_25;
    wire token_15_25;
    wire dep_chan_vld_16_25;
    wire [39:0] dep_chan_data_16_25;
    wire token_16_25;
    wire dep_chan_vld_17_25;
    wire [39:0] dep_chan_data_17_25;
    wire token_17_25;
    wire dep_chan_vld_18_25;
    wire [39:0] dep_chan_data_18_25;
    wire token_18_25;
    wire dep_chan_vld_19_25;
    wire [39:0] dep_chan_data_19_25;
    wire token_19_25;
    wire dep_chan_vld_20_25;
    wire [39:0] dep_chan_data_20_25;
    wire token_20_25;
    wire dep_chan_vld_21_25;
    wire [39:0] dep_chan_data_21_25;
    wire token_21_25;
    wire dep_chan_vld_22_25;
    wire [39:0] dep_chan_data_22_25;
    wire token_22_25;
    wire dep_chan_vld_23_25;
    wire [39:0] dep_chan_data_23_25;
    wire token_23_25;
    wire dep_chan_vld_24_25;
    wire [39:0] dep_chan_data_24_25;
    wire token_24_25;
    wire dep_chan_vld_26_25;
    wire [39:0] dep_chan_data_26_25;
    wire token_26_25;
    wire dep_chan_vld_27_25;
    wire [39:0] dep_chan_data_27_25;
    wire token_27_25;
    wire dep_chan_vld_28_25;
    wire [39:0] dep_chan_data_28_25;
    wire token_28_25;
    wire dep_chan_vld_29_25;
    wire [39:0] dep_chan_data_29_25;
    wire token_29_25;
    wire dep_chan_vld_30_25;
    wire [39:0] dep_chan_data_30_25;
    wire token_30_25;
    wire dep_chan_vld_31_25;
    wire [39:0] dep_chan_data_31_25;
    wire token_31_25;
    wire dep_chan_vld_32_25;
    wire [39:0] dep_chan_data_32_25;
    wire token_32_25;
    wire dep_chan_vld_33_25;
    wire [39:0] dep_chan_data_33_25;
    wire token_33_25;
    wire dep_chan_vld_34_25;
    wire [39:0] dep_chan_data_34_25;
    wire token_34_25;
    wire dep_chan_vld_35_25;
    wire [39:0] dep_chan_data_35_25;
    wire token_35_25;
    wire dep_chan_vld_36_25;
    wire [39:0] dep_chan_data_36_25;
    wire token_36_25;
    wire [32:0] proc_26_data_FIFO_blk;
    wire [32:0] proc_26_data_PIPO_blk;
    wire [32:0] proc_26_start_FIFO_blk;
    wire [32:0] proc_26_TLF_FIFO_blk;
    wire [32:0] proc_26_input_sync_blk;
    wire [32:0] proc_26_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_26;
    reg [32:0] proc_dep_vld_vec_26_reg;
    wire [32:0] in_chan_dep_vld_vec_26;
    wire [1319:0] in_chan_dep_data_vec_26;
    wire [32:0] token_in_vec_26;
    wire [32:0] out_chan_dep_vld_vec_26;
    wire [39:0] out_chan_dep_data_26;
    wire [32:0] token_out_vec_26;
    wire dl_detect_out_26;
    wire dep_chan_vld_0_26;
    wire [39:0] dep_chan_data_0_26;
    wire token_0_26;
    wire dep_chan_vld_1_26;
    wire [39:0] dep_chan_data_1_26;
    wire token_1_26;
    wire dep_chan_vld_3_26;
    wire [39:0] dep_chan_data_3_26;
    wire token_3_26;
    wire dep_chan_vld_6_26;
    wire [39:0] dep_chan_data_6_26;
    wire token_6_26;
    wire dep_chan_vld_7_26;
    wire [39:0] dep_chan_data_7_26;
    wire token_7_26;
    wire dep_chan_vld_8_26;
    wire [39:0] dep_chan_data_8_26;
    wire token_8_26;
    wire dep_chan_vld_9_26;
    wire [39:0] dep_chan_data_9_26;
    wire token_9_26;
    wire dep_chan_vld_10_26;
    wire [39:0] dep_chan_data_10_26;
    wire token_10_26;
    wire dep_chan_vld_11_26;
    wire [39:0] dep_chan_data_11_26;
    wire token_11_26;
    wire dep_chan_vld_12_26;
    wire [39:0] dep_chan_data_12_26;
    wire token_12_26;
    wire dep_chan_vld_13_26;
    wire [39:0] dep_chan_data_13_26;
    wire token_13_26;
    wire dep_chan_vld_14_26;
    wire [39:0] dep_chan_data_14_26;
    wire token_14_26;
    wire dep_chan_vld_15_26;
    wire [39:0] dep_chan_data_15_26;
    wire token_15_26;
    wire dep_chan_vld_16_26;
    wire [39:0] dep_chan_data_16_26;
    wire token_16_26;
    wire dep_chan_vld_17_26;
    wire [39:0] dep_chan_data_17_26;
    wire token_17_26;
    wire dep_chan_vld_18_26;
    wire [39:0] dep_chan_data_18_26;
    wire token_18_26;
    wire dep_chan_vld_19_26;
    wire [39:0] dep_chan_data_19_26;
    wire token_19_26;
    wire dep_chan_vld_20_26;
    wire [39:0] dep_chan_data_20_26;
    wire token_20_26;
    wire dep_chan_vld_21_26;
    wire [39:0] dep_chan_data_21_26;
    wire token_21_26;
    wire dep_chan_vld_22_26;
    wire [39:0] dep_chan_data_22_26;
    wire token_22_26;
    wire dep_chan_vld_23_26;
    wire [39:0] dep_chan_data_23_26;
    wire token_23_26;
    wire dep_chan_vld_24_26;
    wire [39:0] dep_chan_data_24_26;
    wire token_24_26;
    wire dep_chan_vld_25_26;
    wire [39:0] dep_chan_data_25_26;
    wire token_25_26;
    wire dep_chan_vld_27_26;
    wire [39:0] dep_chan_data_27_26;
    wire token_27_26;
    wire dep_chan_vld_28_26;
    wire [39:0] dep_chan_data_28_26;
    wire token_28_26;
    wire dep_chan_vld_29_26;
    wire [39:0] dep_chan_data_29_26;
    wire token_29_26;
    wire dep_chan_vld_30_26;
    wire [39:0] dep_chan_data_30_26;
    wire token_30_26;
    wire dep_chan_vld_31_26;
    wire [39:0] dep_chan_data_31_26;
    wire token_31_26;
    wire dep_chan_vld_32_26;
    wire [39:0] dep_chan_data_32_26;
    wire token_32_26;
    wire dep_chan_vld_33_26;
    wire [39:0] dep_chan_data_33_26;
    wire token_33_26;
    wire dep_chan_vld_34_26;
    wire [39:0] dep_chan_data_34_26;
    wire token_34_26;
    wire dep_chan_vld_35_26;
    wire [39:0] dep_chan_data_35_26;
    wire token_35_26;
    wire dep_chan_vld_36_26;
    wire [39:0] dep_chan_data_36_26;
    wire token_36_26;
    wire [32:0] proc_27_data_FIFO_blk;
    wire [32:0] proc_27_data_PIPO_blk;
    wire [32:0] proc_27_start_FIFO_blk;
    wire [32:0] proc_27_TLF_FIFO_blk;
    wire [32:0] proc_27_input_sync_blk;
    wire [32:0] proc_27_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_27;
    reg [32:0] proc_dep_vld_vec_27_reg;
    wire [32:0] in_chan_dep_vld_vec_27;
    wire [1319:0] in_chan_dep_data_vec_27;
    wire [32:0] token_in_vec_27;
    wire [32:0] out_chan_dep_vld_vec_27;
    wire [39:0] out_chan_dep_data_27;
    wire [32:0] token_out_vec_27;
    wire dl_detect_out_27;
    wire dep_chan_vld_0_27;
    wire [39:0] dep_chan_data_0_27;
    wire token_0_27;
    wire dep_chan_vld_1_27;
    wire [39:0] dep_chan_data_1_27;
    wire token_1_27;
    wire dep_chan_vld_3_27;
    wire [39:0] dep_chan_data_3_27;
    wire token_3_27;
    wire dep_chan_vld_6_27;
    wire [39:0] dep_chan_data_6_27;
    wire token_6_27;
    wire dep_chan_vld_7_27;
    wire [39:0] dep_chan_data_7_27;
    wire token_7_27;
    wire dep_chan_vld_8_27;
    wire [39:0] dep_chan_data_8_27;
    wire token_8_27;
    wire dep_chan_vld_9_27;
    wire [39:0] dep_chan_data_9_27;
    wire token_9_27;
    wire dep_chan_vld_10_27;
    wire [39:0] dep_chan_data_10_27;
    wire token_10_27;
    wire dep_chan_vld_11_27;
    wire [39:0] dep_chan_data_11_27;
    wire token_11_27;
    wire dep_chan_vld_12_27;
    wire [39:0] dep_chan_data_12_27;
    wire token_12_27;
    wire dep_chan_vld_13_27;
    wire [39:0] dep_chan_data_13_27;
    wire token_13_27;
    wire dep_chan_vld_14_27;
    wire [39:0] dep_chan_data_14_27;
    wire token_14_27;
    wire dep_chan_vld_15_27;
    wire [39:0] dep_chan_data_15_27;
    wire token_15_27;
    wire dep_chan_vld_16_27;
    wire [39:0] dep_chan_data_16_27;
    wire token_16_27;
    wire dep_chan_vld_17_27;
    wire [39:0] dep_chan_data_17_27;
    wire token_17_27;
    wire dep_chan_vld_18_27;
    wire [39:0] dep_chan_data_18_27;
    wire token_18_27;
    wire dep_chan_vld_19_27;
    wire [39:0] dep_chan_data_19_27;
    wire token_19_27;
    wire dep_chan_vld_20_27;
    wire [39:0] dep_chan_data_20_27;
    wire token_20_27;
    wire dep_chan_vld_21_27;
    wire [39:0] dep_chan_data_21_27;
    wire token_21_27;
    wire dep_chan_vld_22_27;
    wire [39:0] dep_chan_data_22_27;
    wire token_22_27;
    wire dep_chan_vld_23_27;
    wire [39:0] dep_chan_data_23_27;
    wire token_23_27;
    wire dep_chan_vld_24_27;
    wire [39:0] dep_chan_data_24_27;
    wire token_24_27;
    wire dep_chan_vld_25_27;
    wire [39:0] dep_chan_data_25_27;
    wire token_25_27;
    wire dep_chan_vld_26_27;
    wire [39:0] dep_chan_data_26_27;
    wire token_26_27;
    wire dep_chan_vld_28_27;
    wire [39:0] dep_chan_data_28_27;
    wire token_28_27;
    wire dep_chan_vld_29_27;
    wire [39:0] dep_chan_data_29_27;
    wire token_29_27;
    wire dep_chan_vld_30_27;
    wire [39:0] dep_chan_data_30_27;
    wire token_30_27;
    wire dep_chan_vld_31_27;
    wire [39:0] dep_chan_data_31_27;
    wire token_31_27;
    wire dep_chan_vld_32_27;
    wire [39:0] dep_chan_data_32_27;
    wire token_32_27;
    wire dep_chan_vld_33_27;
    wire [39:0] dep_chan_data_33_27;
    wire token_33_27;
    wire dep_chan_vld_34_27;
    wire [39:0] dep_chan_data_34_27;
    wire token_34_27;
    wire dep_chan_vld_35_27;
    wire [39:0] dep_chan_data_35_27;
    wire token_35_27;
    wire dep_chan_vld_36_27;
    wire [39:0] dep_chan_data_36_27;
    wire token_36_27;
    wire [32:0] proc_28_data_FIFO_blk;
    wire [32:0] proc_28_data_PIPO_blk;
    wire [32:0] proc_28_start_FIFO_blk;
    wire [32:0] proc_28_TLF_FIFO_blk;
    wire [32:0] proc_28_input_sync_blk;
    wire [32:0] proc_28_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_28;
    reg [32:0] proc_dep_vld_vec_28_reg;
    wire [32:0] in_chan_dep_vld_vec_28;
    wire [1319:0] in_chan_dep_data_vec_28;
    wire [32:0] token_in_vec_28;
    wire [32:0] out_chan_dep_vld_vec_28;
    wire [39:0] out_chan_dep_data_28;
    wire [32:0] token_out_vec_28;
    wire dl_detect_out_28;
    wire dep_chan_vld_0_28;
    wire [39:0] dep_chan_data_0_28;
    wire token_0_28;
    wire dep_chan_vld_1_28;
    wire [39:0] dep_chan_data_1_28;
    wire token_1_28;
    wire dep_chan_vld_3_28;
    wire [39:0] dep_chan_data_3_28;
    wire token_3_28;
    wire dep_chan_vld_6_28;
    wire [39:0] dep_chan_data_6_28;
    wire token_6_28;
    wire dep_chan_vld_7_28;
    wire [39:0] dep_chan_data_7_28;
    wire token_7_28;
    wire dep_chan_vld_8_28;
    wire [39:0] dep_chan_data_8_28;
    wire token_8_28;
    wire dep_chan_vld_9_28;
    wire [39:0] dep_chan_data_9_28;
    wire token_9_28;
    wire dep_chan_vld_10_28;
    wire [39:0] dep_chan_data_10_28;
    wire token_10_28;
    wire dep_chan_vld_11_28;
    wire [39:0] dep_chan_data_11_28;
    wire token_11_28;
    wire dep_chan_vld_12_28;
    wire [39:0] dep_chan_data_12_28;
    wire token_12_28;
    wire dep_chan_vld_13_28;
    wire [39:0] dep_chan_data_13_28;
    wire token_13_28;
    wire dep_chan_vld_14_28;
    wire [39:0] dep_chan_data_14_28;
    wire token_14_28;
    wire dep_chan_vld_15_28;
    wire [39:0] dep_chan_data_15_28;
    wire token_15_28;
    wire dep_chan_vld_16_28;
    wire [39:0] dep_chan_data_16_28;
    wire token_16_28;
    wire dep_chan_vld_17_28;
    wire [39:0] dep_chan_data_17_28;
    wire token_17_28;
    wire dep_chan_vld_18_28;
    wire [39:0] dep_chan_data_18_28;
    wire token_18_28;
    wire dep_chan_vld_19_28;
    wire [39:0] dep_chan_data_19_28;
    wire token_19_28;
    wire dep_chan_vld_20_28;
    wire [39:0] dep_chan_data_20_28;
    wire token_20_28;
    wire dep_chan_vld_21_28;
    wire [39:0] dep_chan_data_21_28;
    wire token_21_28;
    wire dep_chan_vld_22_28;
    wire [39:0] dep_chan_data_22_28;
    wire token_22_28;
    wire dep_chan_vld_23_28;
    wire [39:0] dep_chan_data_23_28;
    wire token_23_28;
    wire dep_chan_vld_24_28;
    wire [39:0] dep_chan_data_24_28;
    wire token_24_28;
    wire dep_chan_vld_25_28;
    wire [39:0] dep_chan_data_25_28;
    wire token_25_28;
    wire dep_chan_vld_26_28;
    wire [39:0] dep_chan_data_26_28;
    wire token_26_28;
    wire dep_chan_vld_27_28;
    wire [39:0] dep_chan_data_27_28;
    wire token_27_28;
    wire dep_chan_vld_29_28;
    wire [39:0] dep_chan_data_29_28;
    wire token_29_28;
    wire dep_chan_vld_30_28;
    wire [39:0] dep_chan_data_30_28;
    wire token_30_28;
    wire dep_chan_vld_31_28;
    wire [39:0] dep_chan_data_31_28;
    wire token_31_28;
    wire dep_chan_vld_32_28;
    wire [39:0] dep_chan_data_32_28;
    wire token_32_28;
    wire dep_chan_vld_33_28;
    wire [39:0] dep_chan_data_33_28;
    wire token_33_28;
    wire dep_chan_vld_34_28;
    wire [39:0] dep_chan_data_34_28;
    wire token_34_28;
    wire dep_chan_vld_35_28;
    wire [39:0] dep_chan_data_35_28;
    wire token_35_28;
    wire dep_chan_vld_36_28;
    wire [39:0] dep_chan_data_36_28;
    wire token_36_28;
    wire [32:0] proc_29_data_FIFO_blk;
    wire [32:0] proc_29_data_PIPO_blk;
    wire [32:0] proc_29_start_FIFO_blk;
    wire [32:0] proc_29_TLF_FIFO_blk;
    wire [32:0] proc_29_input_sync_blk;
    wire [32:0] proc_29_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_29;
    reg [32:0] proc_dep_vld_vec_29_reg;
    wire [32:0] in_chan_dep_vld_vec_29;
    wire [1319:0] in_chan_dep_data_vec_29;
    wire [32:0] token_in_vec_29;
    wire [32:0] out_chan_dep_vld_vec_29;
    wire [39:0] out_chan_dep_data_29;
    wire [32:0] token_out_vec_29;
    wire dl_detect_out_29;
    wire dep_chan_vld_0_29;
    wire [39:0] dep_chan_data_0_29;
    wire token_0_29;
    wire dep_chan_vld_1_29;
    wire [39:0] dep_chan_data_1_29;
    wire token_1_29;
    wire dep_chan_vld_3_29;
    wire [39:0] dep_chan_data_3_29;
    wire token_3_29;
    wire dep_chan_vld_6_29;
    wire [39:0] dep_chan_data_6_29;
    wire token_6_29;
    wire dep_chan_vld_7_29;
    wire [39:0] dep_chan_data_7_29;
    wire token_7_29;
    wire dep_chan_vld_8_29;
    wire [39:0] dep_chan_data_8_29;
    wire token_8_29;
    wire dep_chan_vld_9_29;
    wire [39:0] dep_chan_data_9_29;
    wire token_9_29;
    wire dep_chan_vld_10_29;
    wire [39:0] dep_chan_data_10_29;
    wire token_10_29;
    wire dep_chan_vld_11_29;
    wire [39:0] dep_chan_data_11_29;
    wire token_11_29;
    wire dep_chan_vld_12_29;
    wire [39:0] dep_chan_data_12_29;
    wire token_12_29;
    wire dep_chan_vld_13_29;
    wire [39:0] dep_chan_data_13_29;
    wire token_13_29;
    wire dep_chan_vld_14_29;
    wire [39:0] dep_chan_data_14_29;
    wire token_14_29;
    wire dep_chan_vld_15_29;
    wire [39:0] dep_chan_data_15_29;
    wire token_15_29;
    wire dep_chan_vld_16_29;
    wire [39:0] dep_chan_data_16_29;
    wire token_16_29;
    wire dep_chan_vld_17_29;
    wire [39:0] dep_chan_data_17_29;
    wire token_17_29;
    wire dep_chan_vld_18_29;
    wire [39:0] dep_chan_data_18_29;
    wire token_18_29;
    wire dep_chan_vld_19_29;
    wire [39:0] dep_chan_data_19_29;
    wire token_19_29;
    wire dep_chan_vld_20_29;
    wire [39:0] dep_chan_data_20_29;
    wire token_20_29;
    wire dep_chan_vld_21_29;
    wire [39:0] dep_chan_data_21_29;
    wire token_21_29;
    wire dep_chan_vld_22_29;
    wire [39:0] dep_chan_data_22_29;
    wire token_22_29;
    wire dep_chan_vld_23_29;
    wire [39:0] dep_chan_data_23_29;
    wire token_23_29;
    wire dep_chan_vld_24_29;
    wire [39:0] dep_chan_data_24_29;
    wire token_24_29;
    wire dep_chan_vld_25_29;
    wire [39:0] dep_chan_data_25_29;
    wire token_25_29;
    wire dep_chan_vld_26_29;
    wire [39:0] dep_chan_data_26_29;
    wire token_26_29;
    wire dep_chan_vld_27_29;
    wire [39:0] dep_chan_data_27_29;
    wire token_27_29;
    wire dep_chan_vld_28_29;
    wire [39:0] dep_chan_data_28_29;
    wire token_28_29;
    wire dep_chan_vld_30_29;
    wire [39:0] dep_chan_data_30_29;
    wire token_30_29;
    wire dep_chan_vld_31_29;
    wire [39:0] dep_chan_data_31_29;
    wire token_31_29;
    wire dep_chan_vld_32_29;
    wire [39:0] dep_chan_data_32_29;
    wire token_32_29;
    wire dep_chan_vld_33_29;
    wire [39:0] dep_chan_data_33_29;
    wire token_33_29;
    wire dep_chan_vld_34_29;
    wire [39:0] dep_chan_data_34_29;
    wire token_34_29;
    wire dep_chan_vld_35_29;
    wire [39:0] dep_chan_data_35_29;
    wire token_35_29;
    wire dep_chan_vld_36_29;
    wire [39:0] dep_chan_data_36_29;
    wire token_36_29;
    wire [32:0] proc_30_data_FIFO_blk;
    wire [32:0] proc_30_data_PIPO_blk;
    wire [32:0] proc_30_start_FIFO_blk;
    wire [32:0] proc_30_TLF_FIFO_blk;
    wire [32:0] proc_30_input_sync_blk;
    wire [32:0] proc_30_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_30;
    reg [32:0] proc_dep_vld_vec_30_reg;
    wire [32:0] in_chan_dep_vld_vec_30;
    wire [1319:0] in_chan_dep_data_vec_30;
    wire [32:0] token_in_vec_30;
    wire [32:0] out_chan_dep_vld_vec_30;
    wire [39:0] out_chan_dep_data_30;
    wire [32:0] token_out_vec_30;
    wire dl_detect_out_30;
    wire dep_chan_vld_0_30;
    wire [39:0] dep_chan_data_0_30;
    wire token_0_30;
    wire dep_chan_vld_1_30;
    wire [39:0] dep_chan_data_1_30;
    wire token_1_30;
    wire dep_chan_vld_3_30;
    wire [39:0] dep_chan_data_3_30;
    wire token_3_30;
    wire dep_chan_vld_6_30;
    wire [39:0] dep_chan_data_6_30;
    wire token_6_30;
    wire dep_chan_vld_7_30;
    wire [39:0] dep_chan_data_7_30;
    wire token_7_30;
    wire dep_chan_vld_8_30;
    wire [39:0] dep_chan_data_8_30;
    wire token_8_30;
    wire dep_chan_vld_9_30;
    wire [39:0] dep_chan_data_9_30;
    wire token_9_30;
    wire dep_chan_vld_10_30;
    wire [39:0] dep_chan_data_10_30;
    wire token_10_30;
    wire dep_chan_vld_11_30;
    wire [39:0] dep_chan_data_11_30;
    wire token_11_30;
    wire dep_chan_vld_12_30;
    wire [39:0] dep_chan_data_12_30;
    wire token_12_30;
    wire dep_chan_vld_13_30;
    wire [39:0] dep_chan_data_13_30;
    wire token_13_30;
    wire dep_chan_vld_14_30;
    wire [39:0] dep_chan_data_14_30;
    wire token_14_30;
    wire dep_chan_vld_15_30;
    wire [39:0] dep_chan_data_15_30;
    wire token_15_30;
    wire dep_chan_vld_16_30;
    wire [39:0] dep_chan_data_16_30;
    wire token_16_30;
    wire dep_chan_vld_17_30;
    wire [39:0] dep_chan_data_17_30;
    wire token_17_30;
    wire dep_chan_vld_18_30;
    wire [39:0] dep_chan_data_18_30;
    wire token_18_30;
    wire dep_chan_vld_19_30;
    wire [39:0] dep_chan_data_19_30;
    wire token_19_30;
    wire dep_chan_vld_20_30;
    wire [39:0] dep_chan_data_20_30;
    wire token_20_30;
    wire dep_chan_vld_21_30;
    wire [39:0] dep_chan_data_21_30;
    wire token_21_30;
    wire dep_chan_vld_22_30;
    wire [39:0] dep_chan_data_22_30;
    wire token_22_30;
    wire dep_chan_vld_23_30;
    wire [39:0] dep_chan_data_23_30;
    wire token_23_30;
    wire dep_chan_vld_24_30;
    wire [39:0] dep_chan_data_24_30;
    wire token_24_30;
    wire dep_chan_vld_25_30;
    wire [39:0] dep_chan_data_25_30;
    wire token_25_30;
    wire dep_chan_vld_26_30;
    wire [39:0] dep_chan_data_26_30;
    wire token_26_30;
    wire dep_chan_vld_27_30;
    wire [39:0] dep_chan_data_27_30;
    wire token_27_30;
    wire dep_chan_vld_28_30;
    wire [39:0] dep_chan_data_28_30;
    wire token_28_30;
    wire dep_chan_vld_29_30;
    wire [39:0] dep_chan_data_29_30;
    wire token_29_30;
    wire dep_chan_vld_31_30;
    wire [39:0] dep_chan_data_31_30;
    wire token_31_30;
    wire dep_chan_vld_32_30;
    wire [39:0] dep_chan_data_32_30;
    wire token_32_30;
    wire dep_chan_vld_33_30;
    wire [39:0] dep_chan_data_33_30;
    wire token_33_30;
    wire dep_chan_vld_34_30;
    wire [39:0] dep_chan_data_34_30;
    wire token_34_30;
    wire dep_chan_vld_35_30;
    wire [39:0] dep_chan_data_35_30;
    wire token_35_30;
    wire dep_chan_vld_36_30;
    wire [39:0] dep_chan_data_36_30;
    wire token_36_30;
    wire [32:0] proc_31_data_FIFO_blk;
    wire [32:0] proc_31_data_PIPO_blk;
    wire [32:0] proc_31_start_FIFO_blk;
    wire [32:0] proc_31_TLF_FIFO_blk;
    wire [32:0] proc_31_input_sync_blk;
    wire [32:0] proc_31_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_31;
    reg [32:0] proc_dep_vld_vec_31_reg;
    wire [32:0] in_chan_dep_vld_vec_31;
    wire [1319:0] in_chan_dep_data_vec_31;
    wire [32:0] token_in_vec_31;
    wire [32:0] out_chan_dep_vld_vec_31;
    wire [39:0] out_chan_dep_data_31;
    wire [32:0] token_out_vec_31;
    wire dl_detect_out_31;
    wire dep_chan_vld_0_31;
    wire [39:0] dep_chan_data_0_31;
    wire token_0_31;
    wire dep_chan_vld_1_31;
    wire [39:0] dep_chan_data_1_31;
    wire token_1_31;
    wire dep_chan_vld_3_31;
    wire [39:0] dep_chan_data_3_31;
    wire token_3_31;
    wire dep_chan_vld_6_31;
    wire [39:0] dep_chan_data_6_31;
    wire token_6_31;
    wire dep_chan_vld_7_31;
    wire [39:0] dep_chan_data_7_31;
    wire token_7_31;
    wire dep_chan_vld_8_31;
    wire [39:0] dep_chan_data_8_31;
    wire token_8_31;
    wire dep_chan_vld_9_31;
    wire [39:0] dep_chan_data_9_31;
    wire token_9_31;
    wire dep_chan_vld_10_31;
    wire [39:0] dep_chan_data_10_31;
    wire token_10_31;
    wire dep_chan_vld_11_31;
    wire [39:0] dep_chan_data_11_31;
    wire token_11_31;
    wire dep_chan_vld_12_31;
    wire [39:0] dep_chan_data_12_31;
    wire token_12_31;
    wire dep_chan_vld_13_31;
    wire [39:0] dep_chan_data_13_31;
    wire token_13_31;
    wire dep_chan_vld_14_31;
    wire [39:0] dep_chan_data_14_31;
    wire token_14_31;
    wire dep_chan_vld_15_31;
    wire [39:0] dep_chan_data_15_31;
    wire token_15_31;
    wire dep_chan_vld_16_31;
    wire [39:0] dep_chan_data_16_31;
    wire token_16_31;
    wire dep_chan_vld_17_31;
    wire [39:0] dep_chan_data_17_31;
    wire token_17_31;
    wire dep_chan_vld_18_31;
    wire [39:0] dep_chan_data_18_31;
    wire token_18_31;
    wire dep_chan_vld_19_31;
    wire [39:0] dep_chan_data_19_31;
    wire token_19_31;
    wire dep_chan_vld_20_31;
    wire [39:0] dep_chan_data_20_31;
    wire token_20_31;
    wire dep_chan_vld_21_31;
    wire [39:0] dep_chan_data_21_31;
    wire token_21_31;
    wire dep_chan_vld_22_31;
    wire [39:0] dep_chan_data_22_31;
    wire token_22_31;
    wire dep_chan_vld_23_31;
    wire [39:0] dep_chan_data_23_31;
    wire token_23_31;
    wire dep_chan_vld_24_31;
    wire [39:0] dep_chan_data_24_31;
    wire token_24_31;
    wire dep_chan_vld_25_31;
    wire [39:0] dep_chan_data_25_31;
    wire token_25_31;
    wire dep_chan_vld_26_31;
    wire [39:0] dep_chan_data_26_31;
    wire token_26_31;
    wire dep_chan_vld_27_31;
    wire [39:0] dep_chan_data_27_31;
    wire token_27_31;
    wire dep_chan_vld_28_31;
    wire [39:0] dep_chan_data_28_31;
    wire token_28_31;
    wire dep_chan_vld_29_31;
    wire [39:0] dep_chan_data_29_31;
    wire token_29_31;
    wire dep_chan_vld_30_31;
    wire [39:0] dep_chan_data_30_31;
    wire token_30_31;
    wire dep_chan_vld_32_31;
    wire [39:0] dep_chan_data_32_31;
    wire token_32_31;
    wire dep_chan_vld_33_31;
    wire [39:0] dep_chan_data_33_31;
    wire token_33_31;
    wire dep_chan_vld_34_31;
    wire [39:0] dep_chan_data_34_31;
    wire token_34_31;
    wire dep_chan_vld_35_31;
    wire [39:0] dep_chan_data_35_31;
    wire token_35_31;
    wire dep_chan_vld_36_31;
    wire [39:0] dep_chan_data_36_31;
    wire token_36_31;
    wire [32:0] proc_32_data_FIFO_blk;
    wire [32:0] proc_32_data_PIPO_blk;
    wire [32:0] proc_32_start_FIFO_blk;
    wire [32:0] proc_32_TLF_FIFO_blk;
    wire [32:0] proc_32_input_sync_blk;
    wire [32:0] proc_32_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_32;
    reg [32:0] proc_dep_vld_vec_32_reg;
    wire [32:0] in_chan_dep_vld_vec_32;
    wire [1319:0] in_chan_dep_data_vec_32;
    wire [32:0] token_in_vec_32;
    wire [32:0] out_chan_dep_vld_vec_32;
    wire [39:0] out_chan_dep_data_32;
    wire [32:0] token_out_vec_32;
    wire dl_detect_out_32;
    wire dep_chan_vld_0_32;
    wire [39:0] dep_chan_data_0_32;
    wire token_0_32;
    wire dep_chan_vld_1_32;
    wire [39:0] dep_chan_data_1_32;
    wire token_1_32;
    wire dep_chan_vld_3_32;
    wire [39:0] dep_chan_data_3_32;
    wire token_3_32;
    wire dep_chan_vld_6_32;
    wire [39:0] dep_chan_data_6_32;
    wire token_6_32;
    wire dep_chan_vld_7_32;
    wire [39:0] dep_chan_data_7_32;
    wire token_7_32;
    wire dep_chan_vld_8_32;
    wire [39:0] dep_chan_data_8_32;
    wire token_8_32;
    wire dep_chan_vld_9_32;
    wire [39:0] dep_chan_data_9_32;
    wire token_9_32;
    wire dep_chan_vld_10_32;
    wire [39:0] dep_chan_data_10_32;
    wire token_10_32;
    wire dep_chan_vld_11_32;
    wire [39:0] dep_chan_data_11_32;
    wire token_11_32;
    wire dep_chan_vld_12_32;
    wire [39:0] dep_chan_data_12_32;
    wire token_12_32;
    wire dep_chan_vld_13_32;
    wire [39:0] dep_chan_data_13_32;
    wire token_13_32;
    wire dep_chan_vld_14_32;
    wire [39:0] dep_chan_data_14_32;
    wire token_14_32;
    wire dep_chan_vld_15_32;
    wire [39:0] dep_chan_data_15_32;
    wire token_15_32;
    wire dep_chan_vld_16_32;
    wire [39:0] dep_chan_data_16_32;
    wire token_16_32;
    wire dep_chan_vld_17_32;
    wire [39:0] dep_chan_data_17_32;
    wire token_17_32;
    wire dep_chan_vld_18_32;
    wire [39:0] dep_chan_data_18_32;
    wire token_18_32;
    wire dep_chan_vld_19_32;
    wire [39:0] dep_chan_data_19_32;
    wire token_19_32;
    wire dep_chan_vld_20_32;
    wire [39:0] dep_chan_data_20_32;
    wire token_20_32;
    wire dep_chan_vld_21_32;
    wire [39:0] dep_chan_data_21_32;
    wire token_21_32;
    wire dep_chan_vld_22_32;
    wire [39:0] dep_chan_data_22_32;
    wire token_22_32;
    wire dep_chan_vld_23_32;
    wire [39:0] dep_chan_data_23_32;
    wire token_23_32;
    wire dep_chan_vld_24_32;
    wire [39:0] dep_chan_data_24_32;
    wire token_24_32;
    wire dep_chan_vld_25_32;
    wire [39:0] dep_chan_data_25_32;
    wire token_25_32;
    wire dep_chan_vld_26_32;
    wire [39:0] dep_chan_data_26_32;
    wire token_26_32;
    wire dep_chan_vld_27_32;
    wire [39:0] dep_chan_data_27_32;
    wire token_27_32;
    wire dep_chan_vld_28_32;
    wire [39:0] dep_chan_data_28_32;
    wire token_28_32;
    wire dep_chan_vld_29_32;
    wire [39:0] dep_chan_data_29_32;
    wire token_29_32;
    wire dep_chan_vld_30_32;
    wire [39:0] dep_chan_data_30_32;
    wire token_30_32;
    wire dep_chan_vld_31_32;
    wire [39:0] dep_chan_data_31_32;
    wire token_31_32;
    wire dep_chan_vld_33_32;
    wire [39:0] dep_chan_data_33_32;
    wire token_33_32;
    wire dep_chan_vld_34_32;
    wire [39:0] dep_chan_data_34_32;
    wire token_34_32;
    wire dep_chan_vld_35_32;
    wire [39:0] dep_chan_data_35_32;
    wire token_35_32;
    wire dep_chan_vld_36_32;
    wire [39:0] dep_chan_data_36_32;
    wire token_36_32;
    wire [32:0] proc_33_data_FIFO_blk;
    wire [32:0] proc_33_data_PIPO_blk;
    wire [32:0] proc_33_start_FIFO_blk;
    wire [32:0] proc_33_TLF_FIFO_blk;
    wire [32:0] proc_33_input_sync_blk;
    wire [32:0] proc_33_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_33;
    reg [32:0] proc_dep_vld_vec_33_reg;
    wire [32:0] in_chan_dep_vld_vec_33;
    wire [1319:0] in_chan_dep_data_vec_33;
    wire [32:0] token_in_vec_33;
    wire [32:0] out_chan_dep_vld_vec_33;
    wire [39:0] out_chan_dep_data_33;
    wire [32:0] token_out_vec_33;
    wire dl_detect_out_33;
    wire dep_chan_vld_0_33;
    wire [39:0] dep_chan_data_0_33;
    wire token_0_33;
    wire dep_chan_vld_1_33;
    wire [39:0] dep_chan_data_1_33;
    wire token_1_33;
    wire dep_chan_vld_3_33;
    wire [39:0] dep_chan_data_3_33;
    wire token_3_33;
    wire dep_chan_vld_6_33;
    wire [39:0] dep_chan_data_6_33;
    wire token_6_33;
    wire dep_chan_vld_7_33;
    wire [39:0] dep_chan_data_7_33;
    wire token_7_33;
    wire dep_chan_vld_8_33;
    wire [39:0] dep_chan_data_8_33;
    wire token_8_33;
    wire dep_chan_vld_9_33;
    wire [39:0] dep_chan_data_9_33;
    wire token_9_33;
    wire dep_chan_vld_10_33;
    wire [39:0] dep_chan_data_10_33;
    wire token_10_33;
    wire dep_chan_vld_11_33;
    wire [39:0] dep_chan_data_11_33;
    wire token_11_33;
    wire dep_chan_vld_12_33;
    wire [39:0] dep_chan_data_12_33;
    wire token_12_33;
    wire dep_chan_vld_13_33;
    wire [39:0] dep_chan_data_13_33;
    wire token_13_33;
    wire dep_chan_vld_14_33;
    wire [39:0] dep_chan_data_14_33;
    wire token_14_33;
    wire dep_chan_vld_15_33;
    wire [39:0] dep_chan_data_15_33;
    wire token_15_33;
    wire dep_chan_vld_16_33;
    wire [39:0] dep_chan_data_16_33;
    wire token_16_33;
    wire dep_chan_vld_17_33;
    wire [39:0] dep_chan_data_17_33;
    wire token_17_33;
    wire dep_chan_vld_18_33;
    wire [39:0] dep_chan_data_18_33;
    wire token_18_33;
    wire dep_chan_vld_19_33;
    wire [39:0] dep_chan_data_19_33;
    wire token_19_33;
    wire dep_chan_vld_20_33;
    wire [39:0] dep_chan_data_20_33;
    wire token_20_33;
    wire dep_chan_vld_21_33;
    wire [39:0] dep_chan_data_21_33;
    wire token_21_33;
    wire dep_chan_vld_22_33;
    wire [39:0] dep_chan_data_22_33;
    wire token_22_33;
    wire dep_chan_vld_23_33;
    wire [39:0] dep_chan_data_23_33;
    wire token_23_33;
    wire dep_chan_vld_24_33;
    wire [39:0] dep_chan_data_24_33;
    wire token_24_33;
    wire dep_chan_vld_25_33;
    wire [39:0] dep_chan_data_25_33;
    wire token_25_33;
    wire dep_chan_vld_26_33;
    wire [39:0] dep_chan_data_26_33;
    wire token_26_33;
    wire dep_chan_vld_27_33;
    wire [39:0] dep_chan_data_27_33;
    wire token_27_33;
    wire dep_chan_vld_28_33;
    wire [39:0] dep_chan_data_28_33;
    wire token_28_33;
    wire dep_chan_vld_29_33;
    wire [39:0] dep_chan_data_29_33;
    wire token_29_33;
    wire dep_chan_vld_30_33;
    wire [39:0] dep_chan_data_30_33;
    wire token_30_33;
    wire dep_chan_vld_31_33;
    wire [39:0] dep_chan_data_31_33;
    wire token_31_33;
    wire dep_chan_vld_32_33;
    wire [39:0] dep_chan_data_32_33;
    wire token_32_33;
    wire dep_chan_vld_34_33;
    wire [39:0] dep_chan_data_34_33;
    wire token_34_33;
    wire dep_chan_vld_35_33;
    wire [39:0] dep_chan_data_35_33;
    wire token_35_33;
    wire dep_chan_vld_36_33;
    wire [39:0] dep_chan_data_36_33;
    wire token_36_33;
    wire [32:0] proc_34_data_FIFO_blk;
    wire [32:0] proc_34_data_PIPO_blk;
    wire [32:0] proc_34_start_FIFO_blk;
    wire [32:0] proc_34_TLF_FIFO_blk;
    wire [32:0] proc_34_input_sync_blk;
    wire [32:0] proc_34_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_34;
    reg [32:0] proc_dep_vld_vec_34_reg;
    wire [32:0] in_chan_dep_vld_vec_34;
    wire [1319:0] in_chan_dep_data_vec_34;
    wire [32:0] token_in_vec_34;
    wire [32:0] out_chan_dep_vld_vec_34;
    wire [39:0] out_chan_dep_data_34;
    wire [32:0] token_out_vec_34;
    wire dl_detect_out_34;
    wire dep_chan_vld_0_34;
    wire [39:0] dep_chan_data_0_34;
    wire token_0_34;
    wire dep_chan_vld_1_34;
    wire [39:0] dep_chan_data_1_34;
    wire token_1_34;
    wire dep_chan_vld_3_34;
    wire [39:0] dep_chan_data_3_34;
    wire token_3_34;
    wire dep_chan_vld_6_34;
    wire [39:0] dep_chan_data_6_34;
    wire token_6_34;
    wire dep_chan_vld_7_34;
    wire [39:0] dep_chan_data_7_34;
    wire token_7_34;
    wire dep_chan_vld_8_34;
    wire [39:0] dep_chan_data_8_34;
    wire token_8_34;
    wire dep_chan_vld_9_34;
    wire [39:0] dep_chan_data_9_34;
    wire token_9_34;
    wire dep_chan_vld_10_34;
    wire [39:0] dep_chan_data_10_34;
    wire token_10_34;
    wire dep_chan_vld_11_34;
    wire [39:0] dep_chan_data_11_34;
    wire token_11_34;
    wire dep_chan_vld_12_34;
    wire [39:0] dep_chan_data_12_34;
    wire token_12_34;
    wire dep_chan_vld_13_34;
    wire [39:0] dep_chan_data_13_34;
    wire token_13_34;
    wire dep_chan_vld_14_34;
    wire [39:0] dep_chan_data_14_34;
    wire token_14_34;
    wire dep_chan_vld_15_34;
    wire [39:0] dep_chan_data_15_34;
    wire token_15_34;
    wire dep_chan_vld_16_34;
    wire [39:0] dep_chan_data_16_34;
    wire token_16_34;
    wire dep_chan_vld_17_34;
    wire [39:0] dep_chan_data_17_34;
    wire token_17_34;
    wire dep_chan_vld_18_34;
    wire [39:0] dep_chan_data_18_34;
    wire token_18_34;
    wire dep_chan_vld_19_34;
    wire [39:0] dep_chan_data_19_34;
    wire token_19_34;
    wire dep_chan_vld_20_34;
    wire [39:0] dep_chan_data_20_34;
    wire token_20_34;
    wire dep_chan_vld_21_34;
    wire [39:0] dep_chan_data_21_34;
    wire token_21_34;
    wire dep_chan_vld_22_34;
    wire [39:0] dep_chan_data_22_34;
    wire token_22_34;
    wire dep_chan_vld_23_34;
    wire [39:0] dep_chan_data_23_34;
    wire token_23_34;
    wire dep_chan_vld_24_34;
    wire [39:0] dep_chan_data_24_34;
    wire token_24_34;
    wire dep_chan_vld_25_34;
    wire [39:0] dep_chan_data_25_34;
    wire token_25_34;
    wire dep_chan_vld_26_34;
    wire [39:0] dep_chan_data_26_34;
    wire token_26_34;
    wire dep_chan_vld_27_34;
    wire [39:0] dep_chan_data_27_34;
    wire token_27_34;
    wire dep_chan_vld_28_34;
    wire [39:0] dep_chan_data_28_34;
    wire token_28_34;
    wire dep_chan_vld_29_34;
    wire [39:0] dep_chan_data_29_34;
    wire token_29_34;
    wire dep_chan_vld_30_34;
    wire [39:0] dep_chan_data_30_34;
    wire token_30_34;
    wire dep_chan_vld_31_34;
    wire [39:0] dep_chan_data_31_34;
    wire token_31_34;
    wire dep_chan_vld_32_34;
    wire [39:0] dep_chan_data_32_34;
    wire token_32_34;
    wire dep_chan_vld_33_34;
    wire [39:0] dep_chan_data_33_34;
    wire token_33_34;
    wire dep_chan_vld_35_34;
    wire [39:0] dep_chan_data_35_34;
    wire token_35_34;
    wire dep_chan_vld_36_34;
    wire [39:0] dep_chan_data_36_34;
    wire token_36_34;
    wire [32:0] proc_35_data_FIFO_blk;
    wire [32:0] proc_35_data_PIPO_blk;
    wire [32:0] proc_35_start_FIFO_blk;
    wire [32:0] proc_35_TLF_FIFO_blk;
    wire [32:0] proc_35_input_sync_blk;
    wire [32:0] proc_35_output_sync_blk;
    wire [32:0] proc_dep_vld_vec_35;
    reg [32:0] proc_dep_vld_vec_35_reg;
    wire [32:0] in_chan_dep_vld_vec_35;
    wire [1319:0] in_chan_dep_data_vec_35;
    wire [32:0] token_in_vec_35;
    wire [32:0] out_chan_dep_vld_vec_35;
    wire [39:0] out_chan_dep_data_35;
    wire [32:0] token_out_vec_35;
    wire dl_detect_out_35;
    wire dep_chan_vld_0_35;
    wire [39:0] dep_chan_data_0_35;
    wire token_0_35;
    wire dep_chan_vld_1_35;
    wire [39:0] dep_chan_data_1_35;
    wire token_1_35;
    wire dep_chan_vld_3_35;
    wire [39:0] dep_chan_data_3_35;
    wire token_3_35;
    wire dep_chan_vld_6_35;
    wire [39:0] dep_chan_data_6_35;
    wire token_6_35;
    wire dep_chan_vld_7_35;
    wire [39:0] dep_chan_data_7_35;
    wire token_7_35;
    wire dep_chan_vld_8_35;
    wire [39:0] dep_chan_data_8_35;
    wire token_8_35;
    wire dep_chan_vld_9_35;
    wire [39:0] dep_chan_data_9_35;
    wire token_9_35;
    wire dep_chan_vld_10_35;
    wire [39:0] dep_chan_data_10_35;
    wire token_10_35;
    wire dep_chan_vld_11_35;
    wire [39:0] dep_chan_data_11_35;
    wire token_11_35;
    wire dep_chan_vld_12_35;
    wire [39:0] dep_chan_data_12_35;
    wire token_12_35;
    wire dep_chan_vld_13_35;
    wire [39:0] dep_chan_data_13_35;
    wire token_13_35;
    wire dep_chan_vld_14_35;
    wire [39:0] dep_chan_data_14_35;
    wire token_14_35;
    wire dep_chan_vld_15_35;
    wire [39:0] dep_chan_data_15_35;
    wire token_15_35;
    wire dep_chan_vld_16_35;
    wire [39:0] dep_chan_data_16_35;
    wire token_16_35;
    wire dep_chan_vld_17_35;
    wire [39:0] dep_chan_data_17_35;
    wire token_17_35;
    wire dep_chan_vld_18_35;
    wire [39:0] dep_chan_data_18_35;
    wire token_18_35;
    wire dep_chan_vld_19_35;
    wire [39:0] dep_chan_data_19_35;
    wire token_19_35;
    wire dep_chan_vld_20_35;
    wire [39:0] dep_chan_data_20_35;
    wire token_20_35;
    wire dep_chan_vld_21_35;
    wire [39:0] dep_chan_data_21_35;
    wire token_21_35;
    wire dep_chan_vld_22_35;
    wire [39:0] dep_chan_data_22_35;
    wire token_22_35;
    wire dep_chan_vld_23_35;
    wire [39:0] dep_chan_data_23_35;
    wire token_23_35;
    wire dep_chan_vld_24_35;
    wire [39:0] dep_chan_data_24_35;
    wire token_24_35;
    wire dep_chan_vld_25_35;
    wire [39:0] dep_chan_data_25_35;
    wire token_25_35;
    wire dep_chan_vld_26_35;
    wire [39:0] dep_chan_data_26_35;
    wire token_26_35;
    wire dep_chan_vld_27_35;
    wire [39:0] dep_chan_data_27_35;
    wire token_27_35;
    wire dep_chan_vld_28_35;
    wire [39:0] dep_chan_data_28_35;
    wire token_28_35;
    wire dep_chan_vld_29_35;
    wire [39:0] dep_chan_data_29_35;
    wire token_29_35;
    wire dep_chan_vld_30_35;
    wire [39:0] dep_chan_data_30_35;
    wire token_30_35;
    wire dep_chan_vld_31_35;
    wire [39:0] dep_chan_data_31_35;
    wire token_31_35;
    wire dep_chan_vld_32_35;
    wire [39:0] dep_chan_data_32_35;
    wire token_32_35;
    wire dep_chan_vld_33_35;
    wire [39:0] dep_chan_data_33_35;
    wire token_33_35;
    wire dep_chan_vld_34_35;
    wire [39:0] dep_chan_data_34_35;
    wire token_34_35;
    wire dep_chan_vld_36_35;
    wire [39:0] dep_chan_data_36_35;
    wire token_36_35;
    wire [33:0] proc_36_data_FIFO_blk;
    wire [33:0] proc_36_data_PIPO_blk;
    wire [33:0] proc_36_start_FIFO_blk;
    wire [33:0] proc_36_TLF_FIFO_blk;
    wire [33:0] proc_36_input_sync_blk;
    wire [33:0] proc_36_output_sync_blk;
    wire [33:0] proc_dep_vld_vec_36;
    reg [33:0] proc_dep_vld_vec_36_reg;
    wire [33:0] in_chan_dep_vld_vec_36;
    wire [1359:0] in_chan_dep_data_vec_36;
    wire [33:0] token_in_vec_36;
    wire [33:0] out_chan_dep_vld_vec_36;
    wire [39:0] out_chan_dep_data_36;
    wire [33:0] token_out_vec_36;
    wire dl_detect_out_36;
    wire dep_chan_vld_0_36;
    wire [39:0] dep_chan_data_0_36;
    wire token_0_36;
    wire dep_chan_vld_1_36;
    wire [39:0] dep_chan_data_1_36;
    wire token_1_36;
    wire dep_chan_vld_3_36;
    wire [39:0] dep_chan_data_3_36;
    wire token_3_36;
    wire dep_chan_vld_6_36;
    wire [39:0] dep_chan_data_6_36;
    wire token_6_36;
    wire dep_chan_vld_7_36;
    wire [39:0] dep_chan_data_7_36;
    wire token_7_36;
    wire dep_chan_vld_8_36;
    wire [39:0] dep_chan_data_8_36;
    wire token_8_36;
    wire dep_chan_vld_9_36;
    wire [39:0] dep_chan_data_9_36;
    wire token_9_36;
    wire dep_chan_vld_10_36;
    wire [39:0] dep_chan_data_10_36;
    wire token_10_36;
    wire dep_chan_vld_11_36;
    wire [39:0] dep_chan_data_11_36;
    wire token_11_36;
    wire dep_chan_vld_12_36;
    wire [39:0] dep_chan_data_12_36;
    wire token_12_36;
    wire dep_chan_vld_13_36;
    wire [39:0] dep_chan_data_13_36;
    wire token_13_36;
    wire dep_chan_vld_14_36;
    wire [39:0] dep_chan_data_14_36;
    wire token_14_36;
    wire dep_chan_vld_15_36;
    wire [39:0] dep_chan_data_15_36;
    wire token_15_36;
    wire dep_chan_vld_16_36;
    wire [39:0] dep_chan_data_16_36;
    wire token_16_36;
    wire dep_chan_vld_17_36;
    wire [39:0] dep_chan_data_17_36;
    wire token_17_36;
    wire dep_chan_vld_18_36;
    wire [39:0] dep_chan_data_18_36;
    wire token_18_36;
    wire dep_chan_vld_19_36;
    wire [39:0] dep_chan_data_19_36;
    wire token_19_36;
    wire dep_chan_vld_20_36;
    wire [39:0] dep_chan_data_20_36;
    wire token_20_36;
    wire dep_chan_vld_21_36;
    wire [39:0] dep_chan_data_21_36;
    wire token_21_36;
    wire dep_chan_vld_22_36;
    wire [39:0] dep_chan_data_22_36;
    wire token_22_36;
    wire dep_chan_vld_23_36;
    wire [39:0] dep_chan_data_23_36;
    wire token_23_36;
    wire dep_chan_vld_24_36;
    wire [39:0] dep_chan_data_24_36;
    wire token_24_36;
    wire dep_chan_vld_25_36;
    wire [39:0] dep_chan_data_25_36;
    wire token_25_36;
    wire dep_chan_vld_26_36;
    wire [39:0] dep_chan_data_26_36;
    wire token_26_36;
    wire dep_chan_vld_27_36;
    wire [39:0] dep_chan_data_27_36;
    wire token_27_36;
    wire dep_chan_vld_28_36;
    wire [39:0] dep_chan_data_28_36;
    wire token_28_36;
    wire dep_chan_vld_29_36;
    wire [39:0] dep_chan_data_29_36;
    wire token_29_36;
    wire dep_chan_vld_30_36;
    wire [39:0] dep_chan_data_30_36;
    wire token_30_36;
    wire dep_chan_vld_31_36;
    wire [39:0] dep_chan_data_31_36;
    wire token_31_36;
    wire dep_chan_vld_32_36;
    wire [39:0] dep_chan_data_32_36;
    wire token_32_36;
    wire dep_chan_vld_33_36;
    wire [39:0] dep_chan_data_33_36;
    wire token_33_36;
    wire dep_chan_vld_34_36;
    wire [39:0] dep_chan_data_34_36;
    wire token_34_36;
    wire dep_chan_vld_35_36;
    wire [39:0] dep_chan_data_35_36;
    wire token_35_36;
    wire dep_chan_vld_37_36;
    wire [39:0] dep_chan_data_37_36;
    wire token_37_36;
    wire [1:0] proc_37_data_FIFO_blk;
    wire [1:0] proc_37_data_PIPO_blk;
    wire [1:0] proc_37_start_FIFO_blk;
    wire [1:0] proc_37_TLF_FIFO_blk;
    wire [1:0] proc_37_input_sync_blk;
    wire [1:0] proc_37_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_37;
    reg [1:0] proc_dep_vld_vec_37_reg;
    wire [1:0] in_chan_dep_vld_vec_37;
    wire [79:0] in_chan_dep_data_vec_37;
    wire [1:0] token_in_vec_37;
    wire [1:0] out_chan_dep_vld_vec_37;
    wire [39:0] out_chan_dep_data_37;
    wire [1:0] token_out_vec_37;
    wire dl_detect_out_37;
    wire dep_chan_vld_36_37;
    wire [39:0] dep_chan_data_36_37;
    wire token_36_37;
    wire dep_chan_vld_39_37;
    wire [39:0] dep_chan_data_39_37;
    wire token_39_37;
    wire [1:0] proc_38_data_FIFO_blk;
    wire [1:0] proc_38_data_PIPO_blk;
    wire [1:0] proc_38_start_FIFO_blk;
    wire [1:0] proc_38_TLF_FIFO_blk;
    wire [1:0] proc_38_input_sync_blk;
    wire [1:0] proc_38_output_sync_blk;
    wire [1:0] proc_dep_vld_vec_38;
    reg [1:0] proc_dep_vld_vec_38_reg;
    wire [1:0] in_chan_dep_vld_vec_38;
    wire [79:0] in_chan_dep_data_vec_38;
    wire [1:0] token_in_vec_38;
    wire [1:0] out_chan_dep_vld_vec_38;
    wire [39:0] out_chan_dep_data_38;
    wire [1:0] token_out_vec_38;
    wire dl_detect_out_38;
    wire dep_chan_vld_6_38;
    wire [39:0] dep_chan_data_6_38;
    wire token_6_38;
    wire dep_chan_vld_39_38;
    wire [39:0] dep_chan_data_39_38;
    wire token_39_38;
    wire [2:0] proc_39_data_FIFO_blk;
    wire [2:0] proc_39_data_PIPO_blk;
    wire [2:0] proc_39_start_FIFO_blk;
    wire [2:0] proc_39_TLF_FIFO_blk;
    wire [2:0] proc_39_input_sync_blk;
    wire [2:0] proc_39_output_sync_blk;
    wire [2:0] proc_dep_vld_vec_39;
    reg [2:0] proc_dep_vld_vec_39_reg;
    wire [2:0] in_chan_dep_vld_vec_39;
    wire [119:0] in_chan_dep_data_vec_39;
    wire [2:0] token_in_vec_39;
    wire [2:0] out_chan_dep_vld_vec_39;
    wire [39:0] out_chan_dep_data_39;
    wire [2:0] token_out_vec_39;
    wire dl_detect_out_39;
    wire dep_chan_vld_0_39;
    wire [39:0] dep_chan_data_0_39;
    wire token_0_39;
    wire dep_chan_vld_37_39;
    wire [39:0] dep_chan_data_37_39;
    wire token_37_39;
    wire dep_chan_vld_38_39;
    wire [39:0] dep_chan_data_38_39;
    wire token_38_39;
    wire [39:0] dl_in_vec;
    wire dl_detect_out;
    wire token_clear;
    reg [39:0] origin;

    reg ap_done_reg_0;// for module ProcessingElement_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_0 <= 'b0;
        end
        else begin
            ap_done_reg_0 <= ProcessingElement_U0.ap_done & ~ProcessingElement_U0.ap_continue;
        end
    end

    reg ap_done_reg_1;// for module WriteC_U0
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            ap_done_reg_1 <= 'b0;
        end
        else begin
            ap_done_reg_1 <= WriteC_U0.ap_done & ~WriteC_U0.ap_continue;
        end
    end

reg [15:0] trans_in_cnt_0;// for process ReadA_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_0 <= 16'h0;
    end
    else if (ReadA_U0.start_write == 1'b1) begin
        trans_in_cnt_0 <= trans_in_cnt_0 + 16'h1;
    end
    else begin
        trans_in_cnt_0 <= trans_in_cnt_0;
    end
end

reg [15:0] trans_out_cnt_0;// for process ReadA_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_0 <= 16'h0;
    end
    else if (ReadA_U0.ap_done == 1'b1 && ReadA_U0.ap_continue == 1'b1) begin
        trans_out_cnt_0 <= trans_out_cnt_0 + 16'h1;
    end
    else begin
        trans_out_cnt_0 <= trans_out_cnt_0;
    end
end

reg [15:0] trans_in_cnt_1;// for process ReadB_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_1 <= 16'h0;
    end
    else if (ReadB_U0.start_write == 1'b1) begin
        trans_in_cnt_1 <= trans_in_cnt_1 + 16'h1;
    end
    else begin
        trans_in_cnt_1 <= trans_in_cnt_1;
    end
end

reg [15:0] trans_out_cnt_1;// for process ReadB_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_1 <= 16'h0;
    end
    else if (ReadB_U0.ap_done == 1'b1 && ReadB_U0.ap_continue == 1'b1) begin
        trans_out_cnt_1 <= trans_out_cnt_1 + 16'h1;
    end
    else begin
        trans_out_cnt_1 <= trans_out_cnt_1;
    end
end

reg [15:0] trans_in_cnt_2;// for process ConvertWidthB_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_2 <= 16'h0;
    end
    else if (ConvertWidthB_U0.start_write == 1'b1) begin
        trans_in_cnt_2 <= trans_in_cnt_2 + 16'h1;
    end
    else begin
        trans_in_cnt_2 <= trans_in_cnt_2;
    end
end

reg [15:0] trans_out_cnt_2;// for process ConvertWidthB_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_2 <= 16'h0;
    end
    else if (ConvertWidthB_U0.ap_done == 1'b1 && ConvertWidthB_U0.ap_continue == 1'b1) begin
        trans_out_cnt_2 <= trans_out_cnt_2 + 16'h1;
    end
    else begin
        trans_out_cnt_2 <= trans_out_cnt_2;
    end
end

reg [15:0] trans_in_cnt_3;// for process ProcessingElement_31_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_3 <= 16'h0;
    end
    else if (ProcessingElement_31_U0.start_write == 1'b1) begin
        trans_in_cnt_3 <= trans_in_cnt_3 + 16'h1;
    end
    else begin
        trans_in_cnt_3 <= trans_in_cnt_3;
    end
end

reg [15:0] trans_out_cnt_3;// for process ProcessingElement_31_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_3 <= 16'h0;
    end
    else if (ProcessingElement_31_U0.ap_done == 1'b1 && ProcessingElement_31_U0.ap_continue == 1'b1) begin
        trans_out_cnt_3 <= trans_out_cnt_3 + 16'h1;
    end
    else begin
        trans_out_cnt_3 <= trans_out_cnt_3;
    end
end

reg [15:0] trans_in_cnt_4;// for process ProcessingElement_1_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_4 <= 16'h0;
    end
    else if (ProcessingElement_1_U0.start_write == 1'b1) begin
        trans_in_cnt_4 <= trans_in_cnt_4 + 16'h1;
    end
    else begin
        trans_in_cnt_4 <= trans_in_cnt_4;
    end
end

reg [15:0] trans_out_cnt_4;// for process ProcessingElement_1_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_4 <= 16'h0;
    end
    else if (ProcessingElement_1_U0.ap_done == 1'b1 && ProcessingElement_1_U0.ap_continue == 1'b1) begin
        trans_out_cnt_4 <= trans_out_cnt_4 + 16'h1;
    end
    else begin
        trans_out_cnt_4 <= trans_out_cnt_4;
    end
end

reg [15:0] trans_in_cnt_5;// for process entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_in_cnt_5 <= 16'h0;
    end
    else if (entry_proc_U0.start_write == 1'b1) begin
        trans_in_cnt_5 <= trans_in_cnt_5 + 16'h1;
    end
    else begin
        trans_in_cnt_5 <= trans_in_cnt_5;
    end
end

reg [15:0] trans_out_cnt_5;// for process entry_proc_U0
always @(negedge dl_reset or posedge dl_clock) begin
    if (~dl_reset) begin
         trans_out_cnt_5 <= 16'h0;
    end
    else if (entry_proc_U0.ap_done == 1'b1 && entry_proc_U0.ap_continue == 1'b1) begin
        trans_out_cnt_5 <= trans_out_cnt_5 + 16'h1;
    end
    else begin
        trans_out_cnt_5 <= trans_out_cnt_5;
    end
end

    // Process: entry_proc_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 0, 34, 34) MatrixMultiplicationKernel_hls_deadlock_detect_unit_0 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_0),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_0),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_0),
        .token_in_vec(token_in_vec_0),
        .dl_detect_in(dl_detect_out),
        .origin(origin[0]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_0),
        .out_chan_dep_data(out_chan_dep_data_0),
        .token_out_vec(token_out_vec_0),
        .dl_detect_out(dl_in_vec[0]));

    assign proc_0_data_FIFO_blk[0] = 1'b0 | (~entry_proc_U0.c_c_blk_n);
    assign proc_0_data_PIPO_blk[0] = 1'b0;
    assign proc_0_start_FIFO_blk[0] = 1'b0 | (~start_for_WriteC_U0_U.if_full_n & entry_proc_U0.ap_start & ~entry_proc_U0.real_start & (trans_in_cnt_5 == trans_out_cnt_5) & ~start_for_WriteC_U0_U.if_read);
    assign proc_0_TLF_FIFO_blk[0] = 1'b0;
    assign proc_0_input_sync_blk[0] = 1'b0;
    assign proc_0_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_0[0] = dl_detect_out ? proc_dep_vld_vec_0_reg[0] : (proc_0_data_FIFO_blk[0] | proc_0_data_PIPO_blk[0] | proc_0_start_FIFO_blk[0] | proc_0_TLF_FIFO_blk[0] | proc_0_input_sync_blk[0] | proc_0_output_sync_blk[0]);
    assign proc_0_data_FIFO_blk[1] = 1'b0;
    assign proc_0_data_PIPO_blk[1] = 1'b0;
    assign proc_0_start_FIFO_blk[1] = 1'b0;
    assign proc_0_TLF_FIFO_blk[1] = 1'b0;
    assign proc_0_input_sync_blk[1] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_0_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_0[1] = dl_detect_out ? proc_dep_vld_vec_0_reg[1] : (proc_0_data_FIFO_blk[1] | proc_0_data_PIPO_blk[1] | proc_0_start_FIFO_blk[1] | proc_0_TLF_FIFO_blk[1] | proc_0_input_sync_blk[1] | proc_0_output_sync_blk[1]);
    assign proc_0_data_FIFO_blk[2] = 1'b0;
    assign proc_0_data_PIPO_blk[2] = 1'b0;
    assign proc_0_start_FIFO_blk[2] = 1'b0;
    assign proc_0_TLF_FIFO_blk[2] = 1'b0;
    assign proc_0_input_sync_blk[2] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_0_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_0[2] = dl_detect_out ? proc_dep_vld_vec_0_reg[2] : (proc_0_data_FIFO_blk[2] | proc_0_data_PIPO_blk[2] | proc_0_start_FIFO_blk[2] | proc_0_TLF_FIFO_blk[2] | proc_0_input_sync_blk[2] | proc_0_output_sync_blk[2]);
    assign proc_0_data_FIFO_blk[3] = 1'b0;
    assign proc_0_data_PIPO_blk[3] = 1'b0;
    assign proc_0_start_FIFO_blk[3] = 1'b0;
    assign proc_0_TLF_FIFO_blk[3] = 1'b0;
    assign proc_0_input_sync_blk[3] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_0_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_0[3] = dl_detect_out ? proc_dep_vld_vec_0_reg[3] : (proc_0_data_FIFO_blk[3] | proc_0_data_PIPO_blk[3] | proc_0_start_FIFO_blk[3] | proc_0_TLF_FIFO_blk[3] | proc_0_input_sync_blk[3] | proc_0_output_sync_blk[3]);
    assign proc_0_data_FIFO_blk[4] = 1'b0;
    assign proc_0_data_PIPO_blk[4] = 1'b0;
    assign proc_0_start_FIFO_blk[4] = 1'b0;
    assign proc_0_TLF_FIFO_blk[4] = 1'b0;
    assign proc_0_input_sync_blk[4] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_0_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_0[4] = dl_detect_out ? proc_dep_vld_vec_0_reg[4] : (proc_0_data_FIFO_blk[4] | proc_0_data_PIPO_blk[4] | proc_0_start_FIFO_blk[4] | proc_0_TLF_FIFO_blk[4] | proc_0_input_sync_blk[4] | proc_0_output_sync_blk[4]);
    assign proc_0_data_FIFO_blk[5] = 1'b0;
    assign proc_0_data_PIPO_blk[5] = 1'b0;
    assign proc_0_start_FIFO_blk[5] = 1'b0;
    assign proc_0_TLF_FIFO_blk[5] = 1'b0;
    assign proc_0_input_sync_blk[5] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_0_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_0[5] = dl_detect_out ? proc_dep_vld_vec_0_reg[5] : (proc_0_data_FIFO_blk[5] | proc_0_data_PIPO_blk[5] | proc_0_start_FIFO_blk[5] | proc_0_TLF_FIFO_blk[5] | proc_0_input_sync_blk[5] | proc_0_output_sync_blk[5]);
    assign proc_0_data_FIFO_blk[6] = 1'b0;
    assign proc_0_data_PIPO_blk[6] = 1'b0;
    assign proc_0_start_FIFO_blk[6] = 1'b0;
    assign proc_0_TLF_FIFO_blk[6] = 1'b0;
    assign proc_0_input_sync_blk[6] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_0_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_0[6] = dl_detect_out ? proc_dep_vld_vec_0_reg[6] : (proc_0_data_FIFO_blk[6] | proc_0_data_PIPO_blk[6] | proc_0_start_FIFO_blk[6] | proc_0_TLF_FIFO_blk[6] | proc_0_input_sync_blk[6] | proc_0_output_sync_blk[6]);
    assign proc_0_data_FIFO_blk[7] = 1'b0;
    assign proc_0_data_PIPO_blk[7] = 1'b0;
    assign proc_0_start_FIFO_blk[7] = 1'b0;
    assign proc_0_TLF_FIFO_blk[7] = 1'b0;
    assign proc_0_input_sync_blk[7] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_0_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_0[7] = dl_detect_out ? proc_dep_vld_vec_0_reg[7] : (proc_0_data_FIFO_blk[7] | proc_0_data_PIPO_blk[7] | proc_0_start_FIFO_blk[7] | proc_0_TLF_FIFO_blk[7] | proc_0_input_sync_blk[7] | proc_0_output_sync_blk[7]);
    assign proc_0_data_FIFO_blk[8] = 1'b0;
    assign proc_0_data_PIPO_blk[8] = 1'b0;
    assign proc_0_start_FIFO_blk[8] = 1'b0;
    assign proc_0_TLF_FIFO_blk[8] = 1'b0;
    assign proc_0_input_sync_blk[8] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_0_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_0[8] = dl_detect_out ? proc_dep_vld_vec_0_reg[8] : (proc_0_data_FIFO_blk[8] | proc_0_data_PIPO_blk[8] | proc_0_start_FIFO_blk[8] | proc_0_TLF_FIFO_blk[8] | proc_0_input_sync_blk[8] | proc_0_output_sync_blk[8]);
    assign proc_0_data_FIFO_blk[9] = 1'b0;
    assign proc_0_data_PIPO_blk[9] = 1'b0;
    assign proc_0_start_FIFO_blk[9] = 1'b0;
    assign proc_0_TLF_FIFO_blk[9] = 1'b0;
    assign proc_0_input_sync_blk[9] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_0_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_0[9] = dl_detect_out ? proc_dep_vld_vec_0_reg[9] : (proc_0_data_FIFO_blk[9] | proc_0_data_PIPO_blk[9] | proc_0_start_FIFO_blk[9] | proc_0_TLF_FIFO_blk[9] | proc_0_input_sync_blk[9] | proc_0_output_sync_blk[9]);
    assign proc_0_data_FIFO_blk[10] = 1'b0;
    assign proc_0_data_PIPO_blk[10] = 1'b0;
    assign proc_0_start_FIFO_blk[10] = 1'b0;
    assign proc_0_TLF_FIFO_blk[10] = 1'b0;
    assign proc_0_input_sync_blk[10] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_0_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_0[10] = dl_detect_out ? proc_dep_vld_vec_0_reg[10] : (proc_0_data_FIFO_blk[10] | proc_0_data_PIPO_blk[10] | proc_0_start_FIFO_blk[10] | proc_0_TLF_FIFO_blk[10] | proc_0_input_sync_blk[10] | proc_0_output_sync_blk[10]);
    assign proc_0_data_FIFO_blk[11] = 1'b0;
    assign proc_0_data_PIPO_blk[11] = 1'b0;
    assign proc_0_start_FIFO_blk[11] = 1'b0;
    assign proc_0_TLF_FIFO_blk[11] = 1'b0;
    assign proc_0_input_sync_blk[11] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_0_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_0[11] = dl_detect_out ? proc_dep_vld_vec_0_reg[11] : (proc_0_data_FIFO_blk[11] | proc_0_data_PIPO_blk[11] | proc_0_start_FIFO_blk[11] | proc_0_TLF_FIFO_blk[11] | proc_0_input_sync_blk[11] | proc_0_output_sync_blk[11]);
    assign proc_0_data_FIFO_blk[12] = 1'b0;
    assign proc_0_data_PIPO_blk[12] = 1'b0;
    assign proc_0_start_FIFO_blk[12] = 1'b0;
    assign proc_0_TLF_FIFO_blk[12] = 1'b0;
    assign proc_0_input_sync_blk[12] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_0_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_0[12] = dl_detect_out ? proc_dep_vld_vec_0_reg[12] : (proc_0_data_FIFO_blk[12] | proc_0_data_PIPO_blk[12] | proc_0_start_FIFO_blk[12] | proc_0_TLF_FIFO_blk[12] | proc_0_input_sync_blk[12] | proc_0_output_sync_blk[12]);
    assign proc_0_data_FIFO_blk[13] = 1'b0;
    assign proc_0_data_PIPO_blk[13] = 1'b0;
    assign proc_0_start_FIFO_blk[13] = 1'b0;
    assign proc_0_TLF_FIFO_blk[13] = 1'b0;
    assign proc_0_input_sync_blk[13] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_0_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_0[13] = dl_detect_out ? proc_dep_vld_vec_0_reg[13] : (proc_0_data_FIFO_blk[13] | proc_0_data_PIPO_blk[13] | proc_0_start_FIFO_blk[13] | proc_0_TLF_FIFO_blk[13] | proc_0_input_sync_blk[13] | proc_0_output_sync_blk[13]);
    assign proc_0_data_FIFO_blk[14] = 1'b0;
    assign proc_0_data_PIPO_blk[14] = 1'b0;
    assign proc_0_start_FIFO_blk[14] = 1'b0;
    assign proc_0_TLF_FIFO_blk[14] = 1'b0;
    assign proc_0_input_sync_blk[14] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_0_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_0[14] = dl_detect_out ? proc_dep_vld_vec_0_reg[14] : (proc_0_data_FIFO_blk[14] | proc_0_data_PIPO_blk[14] | proc_0_start_FIFO_blk[14] | proc_0_TLF_FIFO_blk[14] | proc_0_input_sync_blk[14] | proc_0_output_sync_blk[14]);
    assign proc_0_data_FIFO_blk[15] = 1'b0;
    assign proc_0_data_PIPO_blk[15] = 1'b0;
    assign proc_0_start_FIFO_blk[15] = 1'b0;
    assign proc_0_TLF_FIFO_blk[15] = 1'b0;
    assign proc_0_input_sync_blk[15] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_0_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_0[15] = dl_detect_out ? proc_dep_vld_vec_0_reg[15] : (proc_0_data_FIFO_blk[15] | proc_0_data_PIPO_blk[15] | proc_0_start_FIFO_blk[15] | proc_0_TLF_FIFO_blk[15] | proc_0_input_sync_blk[15] | proc_0_output_sync_blk[15]);
    assign proc_0_data_FIFO_blk[16] = 1'b0;
    assign proc_0_data_PIPO_blk[16] = 1'b0;
    assign proc_0_start_FIFO_blk[16] = 1'b0;
    assign proc_0_TLF_FIFO_blk[16] = 1'b0;
    assign proc_0_input_sync_blk[16] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_0_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_0[16] = dl_detect_out ? proc_dep_vld_vec_0_reg[16] : (proc_0_data_FIFO_blk[16] | proc_0_data_PIPO_blk[16] | proc_0_start_FIFO_blk[16] | proc_0_TLF_FIFO_blk[16] | proc_0_input_sync_blk[16] | proc_0_output_sync_blk[16]);
    assign proc_0_data_FIFO_blk[17] = 1'b0;
    assign proc_0_data_PIPO_blk[17] = 1'b0;
    assign proc_0_start_FIFO_blk[17] = 1'b0;
    assign proc_0_TLF_FIFO_blk[17] = 1'b0;
    assign proc_0_input_sync_blk[17] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_0_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_0[17] = dl_detect_out ? proc_dep_vld_vec_0_reg[17] : (proc_0_data_FIFO_blk[17] | proc_0_data_PIPO_blk[17] | proc_0_start_FIFO_blk[17] | proc_0_TLF_FIFO_blk[17] | proc_0_input_sync_blk[17] | proc_0_output_sync_blk[17]);
    assign proc_0_data_FIFO_blk[18] = 1'b0;
    assign proc_0_data_PIPO_blk[18] = 1'b0;
    assign proc_0_start_FIFO_blk[18] = 1'b0;
    assign proc_0_TLF_FIFO_blk[18] = 1'b0;
    assign proc_0_input_sync_blk[18] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_0_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_0[18] = dl_detect_out ? proc_dep_vld_vec_0_reg[18] : (proc_0_data_FIFO_blk[18] | proc_0_data_PIPO_blk[18] | proc_0_start_FIFO_blk[18] | proc_0_TLF_FIFO_blk[18] | proc_0_input_sync_blk[18] | proc_0_output_sync_blk[18]);
    assign proc_0_data_FIFO_blk[19] = 1'b0;
    assign proc_0_data_PIPO_blk[19] = 1'b0;
    assign proc_0_start_FIFO_blk[19] = 1'b0;
    assign proc_0_TLF_FIFO_blk[19] = 1'b0;
    assign proc_0_input_sync_blk[19] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_0_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_0[19] = dl_detect_out ? proc_dep_vld_vec_0_reg[19] : (proc_0_data_FIFO_blk[19] | proc_0_data_PIPO_blk[19] | proc_0_start_FIFO_blk[19] | proc_0_TLF_FIFO_blk[19] | proc_0_input_sync_blk[19] | proc_0_output_sync_blk[19]);
    assign proc_0_data_FIFO_blk[20] = 1'b0;
    assign proc_0_data_PIPO_blk[20] = 1'b0;
    assign proc_0_start_FIFO_blk[20] = 1'b0;
    assign proc_0_TLF_FIFO_blk[20] = 1'b0;
    assign proc_0_input_sync_blk[20] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_0_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_0[20] = dl_detect_out ? proc_dep_vld_vec_0_reg[20] : (proc_0_data_FIFO_blk[20] | proc_0_data_PIPO_blk[20] | proc_0_start_FIFO_blk[20] | proc_0_TLF_FIFO_blk[20] | proc_0_input_sync_blk[20] | proc_0_output_sync_blk[20]);
    assign proc_0_data_FIFO_blk[21] = 1'b0;
    assign proc_0_data_PIPO_blk[21] = 1'b0;
    assign proc_0_start_FIFO_blk[21] = 1'b0;
    assign proc_0_TLF_FIFO_blk[21] = 1'b0;
    assign proc_0_input_sync_blk[21] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_0_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_0[21] = dl_detect_out ? proc_dep_vld_vec_0_reg[21] : (proc_0_data_FIFO_blk[21] | proc_0_data_PIPO_blk[21] | proc_0_start_FIFO_blk[21] | proc_0_TLF_FIFO_blk[21] | proc_0_input_sync_blk[21] | proc_0_output_sync_blk[21]);
    assign proc_0_data_FIFO_blk[22] = 1'b0;
    assign proc_0_data_PIPO_blk[22] = 1'b0;
    assign proc_0_start_FIFO_blk[22] = 1'b0;
    assign proc_0_TLF_FIFO_blk[22] = 1'b0;
    assign proc_0_input_sync_blk[22] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_0_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_0[22] = dl_detect_out ? proc_dep_vld_vec_0_reg[22] : (proc_0_data_FIFO_blk[22] | proc_0_data_PIPO_blk[22] | proc_0_start_FIFO_blk[22] | proc_0_TLF_FIFO_blk[22] | proc_0_input_sync_blk[22] | proc_0_output_sync_blk[22]);
    assign proc_0_data_FIFO_blk[23] = 1'b0;
    assign proc_0_data_PIPO_blk[23] = 1'b0;
    assign proc_0_start_FIFO_blk[23] = 1'b0;
    assign proc_0_TLF_FIFO_blk[23] = 1'b0;
    assign proc_0_input_sync_blk[23] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_0_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_0[23] = dl_detect_out ? proc_dep_vld_vec_0_reg[23] : (proc_0_data_FIFO_blk[23] | proc_0_data_PIPO_blk[23] | proc_0_start_FIFO_blk[23] | proc_0_TLF_FIFO_blk[23] | proc_0_input_sync_blk[23] | proc_0_output_sync_blk[23]);
    assign proc_0_data_FIFO_blk[24] = 1'b0;
    assign proc_0_data_PIPO_blk[24] = 1'b0;
    assign proc_0_start_FIFO_blk[24] = 1'b0;
    assign proc_0_TLF_FIFO_blk[24] = 1'b0;
    assign proc_0_input_sync_blk[24] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_0_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_0[24] = dl_detect_out ? proc_dep_vld_vec_0_reg[24] : (proc_0_data_FIFO_blk[24] | proc_0_data_PIPO_blk[24] | proc_0_start_FIFO_blk[24] | proc_0_TLF_FIFO_blk[24] | proc_0_input_sync_blk[24] | proc_0_output_sync_blk[24]);
    assign proc_0_data_FIFO_blk[25] = 1'b0;
    assign proc_0_data_PIPO_blk[25] = 1'b0;
    assign proc_0_start_FIFO_blk[25] = 1'b0;
    assign proc_0_TLF_FIFO_blk[25] = 1'b0;
    assign proc_0_input_sync_blk[25] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_0_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_0[25] = dl_detect_out ? proc_dep_vld_vec_0_reg[25] : (proc_0_data_FIFO_blk[25] | proc_0_data_PIPO_blk[25] | proc_0_start_FIFO_blk[25] | proc_0_TLF_FIFO_blk[25] | proc_0_input_sync_blk[25] | proc_0_output_sync_blk[25]);
    assign proc_0_data_FIFO_blk[26] = 1'b0;
    assign proc_0_data_PIPO_blk[26] = 1'b0;
    assign proc_0_start_FIFO_blk[26] = 1'b0;
    assign proc_0_TLF_FIFO_blk[26] = 1'b0;
    assign proc_0_input_sync_blk[26] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_0_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_0[26] = dl_detect_out ? proc_dep_vld_vec_0_reg[26] : (proc_0_data_FIFO_blk[26] | proc_0_data_PIPO_blk[26] | proc_0_start_FIFO_blk[26] | proc_0_TLF_FIFO_blk[26] | proc_0_input_sync_blk[26] | proc_0_output_sync_blk[26]);
    assign proc_0_data_FIFO_blk[27] = 1'b0;
    assign proc_0_data_PIPO_blk[27] = 1'b0;
    assign proc_0_start_FIFO_blk[27] = 1'b0;
    assign proc_0_TLF_FIFO_blk[27] = 1'b0;
    assign proc_0_input_sync_blk[27] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_0_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_0[27] = dl_detect_out ? proc_dep_vld_vec_0_reg[27] : (proc_0_data_FIFO_blk[27] | proc_0_data_PIPO_blk[27] | proc_0_start_FIFO_blk[27] | proc_0_TLF_FIFO_blk[27] | proc_0_input_sync_blk[27] | proc_0_output_sync_blk[27]);
    assign proc_0_data_FIFO_blk[28] = 1'b0;
    assign proc_0_data_PIPO_blk[28] = 1'b0;
    assign proc_0_start_FIFO_blk[28] = 1'b0;
    assign proc_0_TLF_FIFO_blk[28] = 1'b0;
    assign proc_0_input_sync_blk[28] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_0_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_0[28] = dl_detect_out ? proc_dep_vld_vec_0_reg[28] : (proc_0_data_FIFO_blk[28] | proc_0_data_PIPO_blk[28] | proc_0_start_FIFO_blk[28] | proc_0_TLF_FIFO_blk[28] | proc_0_input_sync_blk[28] | proc_0_output_sync_blk[28]);
    assign proc_0_data_FIFO_blk[29] = 1'b0;
    assign proc_0_data_PIPO_blk[29] = 1'b0;
    assign proc_0_start_FIFO_blk[29] = 1'b0;
    assign proc_0_TLF_FIFO_blk[29] = 1'b0;
    assign proc_0_input_sync_blk[29] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_0_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_0[29] = dl_detect_out ? proc_dep_vld_vec_0_reg[29] : (proc_0_data_FIFO_blk[29] | proc_0_data_PIPO_blk[29] | proc_0_start_FIFO_blk[29] | proc_0_TLF_FIFO_blk[29] | proc_0_input_sync_blk[29] | proc_0_output_sync_blk[29]);
    assign proc_0_data_FIFO_blk[30] = 1'b0;
    assign proc_0_data_PIPO_blk[30] = 1'b0;
    assign proc_0_start_FIFO_blk[30] = 1'b0;
    assign proc_0_TLF_FIFO_blk[30] = 1'b0;
    assign proc_0_input_sync_blk[30] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_0_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_0[30] = dl_detect_out ? proc_dep_vld_vec_0_reg[30] : (proc_0_data_FIFO_blk[30] | proc_0_data_PIPO_blk[30] | proc_0_start_FIFO_blk[30] | proc_0_TLF_FIFO_blk[30] | proc_0_input_sync_blk[30] | proc_0_output_sync_blk[30]);
    assign proc_0_data_FIFO_blk[31] = 1'b0;
    assign proc_0_data_PIPO_blk[31] = 1'b0;
    assign proc_0_start_FIFO_blk[31] = 1'b0;
    assign proc_0_TLF_FIFO_blk[31] = 1'b0;
    assign proc_0_input_sync_blk[31] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_0_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_0[31] = dl_detect_out ? proc_dep_vld_vec_0_reg[31] : (proc_0_data_FIFO_blk[31] | proc_0_data_PIPO_blk[31] | proc_0_start_FIFO_blk[31] | proc_0_TLF_FIFO_blk[31] | proc_0_input_sync_blk[31] | proc_0_output_sync_blk[31]);
    assign proc_0_data_FIFO_blk[32] = 1'b0;
    assign proc_0_data_PIPO_blk[32] = 1'b0;
    assign proc_0_start_FIFO_blk[32] = 1'b0;
    assign proc_0_TLF_FIFO_blk[32] = 1'b0;
    assign proc_0_input_sync_blk[32] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_0_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_0[32] = dl_detect_out ? proc_dep_vld_vec_0_reg[32] : (proc_0_data_FIFO_blk[32] | proc_0_data_PIPO_blk[32] | proc_0_start_FIFO_blk[32] | proc_0_TLF_FIFO_blk[32] | proc_0_input_sync_blk[32] | proc_0_output_sync_blk[32]);
    assign proc_0_data_FIFO_blk[33] = 1'b0;
    assign proc_0_data_PIPO_blk[33] = 1'b0;
    assign proc_0_start_FIFO_blk[33] = 1'b0;
    assign proc_0_TLF_FIFO_blk[33] = 1'b0;
    assign proc_0_input_sync_blk[33] = 1'b0 | (ap_sync_entry_proc_U0_ap_ready & entry_proc_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_0_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_0[33] = dl_detect_out ? proc_dep_vld_vec_0_reg[33] : (proc_0_data_FIFO_blk[33] | proc_0_data_PIPO_blk[33] | proc_0_start_FIFO_blk[33] | proc_0_TLF_FIFO_blk[33] | proc_0_input_sync_blk[33] | proc_0_output_sync_blk[33]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_0_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_0_reg <= proc_dep_vld_vec_0;
        end
    end
    assign in_chan_dep_vld_vec_0[0] = dep_chan_vld_1_0;
    assign in_chan_dep_data_vec_0[39 : 0] = dep_chan_data_1_0;
    assign token_in_vec_0[0] = token_1_0;
    assign in_chan_dep_vld_vec_0[1] = dep_chan_vld_3_0;
    assign in_chan_dep_data_vec_0[79 : 40] = dep_chan_data_3_0;
    assign token_in_vec_0[1] = token_3_0;
    assign in_chan_dep_vld_vec_0[2] = dep_chan_vld_6_0;
    assign in_chan_dep_data_vec_0[119 : 80] = dep_chan_data_6_0;
    assign token_in_vec_0[2] = token_6_0;
    assign in_chan_dep_vld_vec_0[3] = dep_chan_vld_7_0;
    assign in_chan_dep_data_vec_0[159 : 120] = dep_chan_data_7_0;
    assign token_in_vec_0[3] = token_7_0;
    assign in_chan_dep_vld_vec_0[4] = dep_chan_vld_8_0;
    assign in_chan_dep_data_vec_0[199 : 160] = dep_chan_data_8_0;
    assign token_in_vec_0[4] = token_8_0;
    assign in_chan_dep_vld_vec_0[5] = dep_chan_vld_9_0;
    assign in_chan_dep_data_vec_0[239 : 200] = dep_chan_data_9_0;
    assign token_in_vec_0[5] = token_9_0;
    assign in_chan_dep_vld_vec_0[6] = dep_chan_vld_10_0;
    assign in_chan_dep_data_vec_0[279 : 240] = dep_chan_data_10_0;
    assign token_in_vec_0[6] = token_10_0;
    assign in_chan_dep_vld_vec_0[7] = dep_chan_vld_11_0;
    assign in_chan_dep_data_vec_0[319 : 280] = dep_chan_data_11_0;
    assign token_in_vec_0[7] = token_11_0;
    assign in_chan_dep_vld_vec_0[8] = dep_chan_vld_12_0;
    assign in_chan_dep_data_vec_0[359 : 320] = dep_chan_data_12_0;
    assign token_in_vec_0[8] = token_12_0;
    assign in_chan_dep_vld_vec_0[9] = dep_chan_vld_13_0;
    assign in_chan_dep_data_vec_0[399 : 360] = dep_chan_data_13_0;
    assign token_in_vec_0[9] = token_13_0;
    assign in_chan_dep_vld_vec_0[10] = dep_chan_vld_14_0;
    assign in_chan_dep_data_vec_0[439 : 400] = dep_chan_data_14_0;
    assign token_in_vec_0[10] = token_14_0;
    assign in_chan_dep_vld_vec_0[11] = dep_chan_vld_15_0;
    assign in_chan_dep_data_vec_0[479 : 440] = dep_chan_data_15_0;
    assign token_in_vec_0[11] = token_15_0;
    assign in_chan_dep_vld_vec_0[12] = dep_chan_vld_16_0;
    assign in_chan_dep_data_vec_0[519 : 480] = dep_chan_data_16_0;
    assign token_in_vec_0[12] = token_16_0;
    assign in_chan_dep_vld_vec_0[13] = dep_chan_vld_17_0;
    assign in_chan_dep_data_vec_0[559 : 520] = dep_chan_data_17_0;
    assign token_in_vec_0[13] = token_17_0;
    assign in_chan_dep_vld_vec_0[14] = dep_chan_vld_18_0;
    assign in_chan_dep_data_vec_0[599 : 560] = dep_chan_data_18_0;
    assign token_in_vec_0[14] = token_18_0;
    assign in_chan_dep_vld_vec_0[15] = dep_chan_vld_19_0;
    assign in_chan_dep_data_vec_0[639 : 600] = dep_chan_data_19_0;
    assign token_in_vec_0[15] = token_19_0;
    assign in_chan_dep_vld_vec_0[16] = dep_chan_vld_20_0;
    assign in_chan_dep_data_vec_0[679 : 640] = dep_chan_data_20_0;
    assign token_in_vec_0[16] = token_20_0;
    assign in_chan_dep_vld_vec_0[17] = dep_chan_vld_21_0;
    assign in_chan_dep_data_vec_0[719 : 680] = dep_chan_data_21_0;
    assign token_in_vec_0[17] = token_21_0;
    assign in_chan_dep_vld_vec_0[18] = dep_chan_vld_22_0;
    assign in_chan_dep_data_vec_0[759 : 720] = dep_chan_data_22_0;
    assign token_in_vec_0[18] = token_22_0;
    assign in_chan_dep_vld_vec_0[19] = dep_chan_vld_23_0;
    assign in_chan_dep_data_vec_0[799 : 760] = dep_chan_data_23_0;
    assign token_in_vec_0[19] = token_23_0;
    assign in_chan_dep_vld_vec_0[20] = dep_chan_vld_24_0;
    assign in_chan_dep_data_vec_0[839 : 800] = dep_chan_data_24_0;
    assign token_in_vec_0[20] = token_24_0;
    assign in_chan_dep_vld_vec_0[21] = dep_chan_vld_25_0;
    assign in_chan_dep_data_vec_0[879 : 840] = dep_chan_data_25_0;
    assign token_in_vec_0[21] = token_25_0;
    assign in_chan_dep_vld_vec_0[22] = dep_chan_vld_26_0;
    assign in_chan_dep_data_vec_0[919 : 880] = dep_chan_data_26_0;
    assign token_in_vec_0[22] = token_26_0;
    assign in_chan_dep_vld_vec_0[23] = dep_chan_vld_27_0;
    assign in_chan_dep_data_vec_0[959 : 920] = dep_chan_data_27_0;
    assign token_in_vec_0[23] = token_27_0;
    assign in_chan_dep_vld_vec_0[24] = dep_chan_vld_28_0;
    assign in_chan_dep_data_vec_0[999 : 960] = dep_chan_data_28_0;
    assign token_in_vec_0[24] = token_28_0;
    assign in_chan_dep_vld_vec_0[25] = dep_chan_vld_29_0;
    assign in_chan_dep_data_vec_0[1039 : 1000] = dep_chan_data_29_0;
    assign token_in_vec_0[25] = token_29_0;
    assign in_chan_dep_vld_vec_0[26] = dep_chan_vld_30_0;
    assign in_chan_dep_data_vec_0[1079 : 1040] = dep_chan_data_30_0;
    assign token_in_vec_0[26] = token_30_0;
    assign in_chan_dep_vld_vec_0[27] = dep_chan_vld_31_0;
    assign in_chan_dep_data_vec_0[1119 : 1080] = dep_chan_data_31_0;
    assign token_in_vec_0[27] = token_31_0;
    assign in_chan_dep_vld_vec_0[28] = dep_chan_vld_32_0;
    assign in_chan_dep_data_vec_0[1159 : 1120] = dep_chan_data_32_0;
    assign token_in_vec_0[28] = token_32_0;
    assign in_chan_dep_vld_vec_0[29] = dep_chan_vld_33_0;
    assign in_chan_dep_data_vec_0[1199 : 1160] = dep_chan_data_33_0;
    assign token_in_vec_0[29] = token_33_0;
    assign in_chan_dep_vld_vec_0[30] = dep_chan_vld_34_0;
    assign in_chan_dep_data_vec_0[1239 : 1200] = dep_chan_data_34_0;
    assign token_in_vec_0[30] = token_34_0;
    assign in_chan_dep_vld_vec_0[31] = dep_chan_vld_35_0;
    assign in_chan_dep_data_vec_0[1279 : 1240] = dep_chan_data_35_0;
    assign token_in_vec_0[31] = token_35_0;
    assign in_chan_dep_vld_vec_0[32] = dep_chan_vld_36_0;
    assign in_chan_dep_data_vec_0[1319 : 1280] = dep_chan_data_36_0;
    assign token_in_vec_0[32] = token_36_0;
    assign in_chan_dep_vld_vec_0[33] = dep_chan_vld_39_0;
    assign in_chan_dep_data_vec_0[1359 : 1320] = dep_chan_data_39_0;
    assign token_in_vec_0[33] = token_39_0;
    assign dep_chan_vld_0_39 = out_chan_dep_vld_vec_0[0];
    assign dep_chan_data_0_39 = out_chan_dep_data_0;
    assign token_0_39 = token_out_vec_0[0];
    assign dep_chan_vld_0_1 = out_chan_dep_vld_vec_0[1];
    assign dep_chan_data_0_1 = out_chan_dep_data_0;
    assign token_0_1 = token_out_vec_0[1];
    assign dep_chan_vld_0_3 = out_chan_dep_vld_vec_0[2];
    assign dep_chan_data_0_3 = out_chan_dep_data_0;
    assign token_0_3 = token_out_vec_0[2];
    assign dep_chan_vld_0_6 = out_chan_dep_vld_vec_0[3];
    assign dep_chan_data_0_6 = out_chan_dep_data_0;
    assign token_0_6 = token_out_vec_0[3];
    assign dep_chan_vld_0_7 = out_chan_dep_vld_vec_0[4];
    assign dep_chan_data_0_7 = out_chan_dep_data_0;
    assign token_0_7 = token_out_vec_0[4];
    assign dep_chan_vld_0_8 = out_chan_dep_vld_vec_0[5];
    assign dep_chan_data_0_8 = out_chan_dep_data_0;
    assign token_0_8 = token_out_vec_0[5];
    assign dep_chan_vld_0_9 = out_chan_dep_vld_vec_0[6];
    assign dep_chan_data_0_9 = out_chan_dep_data_0;
    assign token_0_9 = token_out_vec_0[6];
    assign dep_chan_vld_0_10 = out_chan_dep_vld_vec_0[7];
    assign dep_chan_data_0_10 = out_chan_dep_data_0;
    assign token_0_10 = token_out_vec_0[7];
    assign dep_chan_vld_0_11 = out_chan_dep_vld_vec_0[8];
    assign dep_chan_data_0_11 = out_chan_dep_data_0;
    assign token_0_11 = token_out_vec_0[8];
    assign dep_chan_vld_0_12 = out_chan_dep_vld_vec_0[9];
    assign dep_chan_data_0_12 = out_chan_dep_data_0;
    assign token_0_12 = token_out_vec_0[9];
    assign dep_chan_vld_0_13 = out_chan_dep_vld_vec_0[10];
    assign dep_chan_data_0_13 = out_chan_dep_data_0;
    assign token_0_13 = token_out_vec_0[10];
    assign dep_chan_vld_0_14 = out_chan_dep_vld_vec_0[11];
    assign dep_chan_data_0_14 = out_chan_dep_data_0;
    assign token_0_14 = token_out_vec_0[11];
    assign dep_chan_vld_0_15 = out_chan_dep_vld_vec_0[12];
    assign dep_chan_data_0_15 = out_chan_dep_data_0;
    assign token_0_15 = token_out_vec_0[12];
    assign dep_chan_vld_0_16 = out_chan_dep_vld_vec_0[13];
    assign dep_chan_data_0_16 = out_chan_dep_data_0;
    assign token_0_16 = token_out_vec_0[13];
    assign dep_chan_vld_0_17 = out_chan_dep_vld_vec_0[14];
    assign dep_chan_data_0_17 = out_chan_dep_data_0;
    assign token_0_17 = token_out_vec_0[14];
    assign dep_chan_vld_0_18 = out_chan_dep_vld_vec_0[15];
    assign dep_chan_data_0_18 = out_chan_dep_data_0;
    assign token_0_18 = token_out_vec_0[15];
    assign dep_chan_vld_0_19 = out_chan_dep_vld_vec_0[16];
    assign dep_chan_data_0_19 = out_chan_dep_data_0;
    assign token_0_19 = token_out_vec_0[16];
    assign dep_chan_vld_0_20 = out_chan_dep_vld_vec_0[17];
    assign dep_chan_data_0_20 = out_chan_dep_data_0;
    assign token_0_20 = token_out_vec_0[17];
    assign dep_chan_vld_0_21 = out_chan_dep_vld_vec_0[18];
    assign dep_chan_data_0_21 = out_chan_dep_data_0;
    assign token_0_21 = token_out_vec_0[18];
    assign dep_chan_vld_0_22 = out_chan_dep_vld_vec_0[19];
    assign dep_chan_data_0_22 = out_chan_dep_data_0;
    assign token_0_22 = token_out_vec_0[19];
    assign dep_chan_vld_0_23 = out_chan_dep_vld_vec_0[20];
    assign dep_chan_data_0_23 = out_chan_dep_data_0;
    assign token_0_23 = token_out_vec_0[20];
    assign dep_chan_vld_0_24 = out_chan_dep_vld_vec_0[21];
    assign dep_chan_data_0_24 = out_chan_dep_data_0;
    assign token_0_24 = token_out_vec_0[21];
    assign dep_chan_vld_0_25 = out_chan_dep_vld_vec_0[22];
    assign dep_chan_data_0_25 = out_chan_dep_data_0;
    assign token_0_25 = token_out_vec_0[22];
    assign dep_chan_vld_0_26 = out_chan_dep_vld_vec_0[23];
    assign dep_chan_data_0_26 = out_chan_dep_data_0;
    assign token_0_26 = token_out_vec_0[23];
    assign dep_chan_vld_0_27 = out_chan_dep_vld_vec_0[24];
    assign dep_chan_data_0_27 = out_chan_dep_data_0;
    assign token_0_27 = token_out_vec_0[24];
    assign dep_chan_vld_0_28 = out_chan_dep_vld_vec_0[25];
    assign dep_chan_data_0_28 = out_chan_dep_data_0;
    assign token_0_28 = token_out_vec_0[25];
    assign dep_chan_vld_0_29 = out_chan_dep_vld_vec_0[26];
    assign dep_chan_data_0_29 = out_chan_dep_data_0;
    assign token_0_29 = token_out_vec_0[26];
    assign dep_chan_vld_0_30 = out_chan_dep_vld_vec_0[27];
    assign dep_chan_data_0_30 = out_chan_dep_data_0;
    assign token_0_30 = token_out_vec_0[27];
    assign dep_chan_vld_0_31 = out_chan_dep_vld_vec_0[28];
    assign dep_chan_data_0_31 = out_chan_dep_data_0;
    assign token_0_31 = token_out_vec_0[28];
    assign dep_chan_vld_0_32 = out_chan_dep_vld_vec_0[29];
    assign dep_chan_data_0_32 = out_chan_dep_data_0;
    assign token_0_32 = token_out_vec_0[29];
    assign dep_chan_vld_0_33 = out_chan_dep_vld_vec_0[30];
    assign dep_chan_data_0_33 = out_chan_dep_data_0;
    assign token_0_33 = token_out_vec_0[30];
    assign dep_chan_vld_0_34 = out_chan_dep_vld_vec_0[31];
    assign dep_chan_data_0_34 = out_chan_dep_data_0;
    assign token_0_34 = token_out_vec_0[31];
    assign dep_chan_vld_0_35 = out_chan_dep_vld_vec_0[32];
    assign dep_chan_data_0_35 = out_chan_dep_data_0;
    assign token_0_35 = token_out_vec_0[32];
    assign dep_chan_vld_0_36 = out_chan_dep_vld_vec_0[33];
    assign dep_chan_data_0_36 = out_chan_dep_data_0;
    assign token_0_36 = token_out_vec_0[33];

    // Process: ReadA_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 1, 34, 34) MatrixMultiplicationKernel_hls_deadlock_detect_unit_1 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_1),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_1),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_1),
        .token_in_vec(token_in_vec_1),
        .dl_detect_in(dl_detect_out),
        .origin(origin[1]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_1),
        .out_chan_dep_data(out_chan_dep_data_1),
        .token_out_vec(token_out_vec_1),
        .dl_detect_out(dl_in_vec[1]));

    assign proc_1_data_FIFO_blk[0] = 1'b0 | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_0_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_1_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_2_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_3_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_4_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_5_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_6_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_7_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_8_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_9_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_10_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_11_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_12_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_13_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_14_blk_n) | (~ReadA_U0.grp_ReadA_Pipeline_ReadA_N0_ReadA_M0_ReadA_K0_ReadA_N1_ReadA_N2_fu_152.aSplit_15_blk_n) | (~ReadA_U0.size_n_c5_blk_n) | (~ReadA_U0.size_k_c8_blk_n) | (~ReadA_U0.size_m_c13_blk_n);
    assign proc_1_data_PIPO_blk[0] = 1'b0;
    assign proc_1_start_FIFO_blk[0] = 1'b0 | (~start_for_TransposeA_U0_U.if_full_n & ReadA_U0.ap_start & ~ReadA_U0.real_start & (trans_in_cnt_0 == trans_out_cnt_0) & ~start_for_TransposeA_U0_U.if_read);
    assign proc_1_TLF_FIFO_blk[0] = 1'b0;
    assign proc_1_input_sync_blk[0] = 1'b0;
    assign proc_1_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_1[0] = dl_detect_out ? proc_dep_vld_vec_1_reg[0] : (proc_1_data_FIFO_blk[0] | proc_1_data_PIPO_blk[0] | proc_1_start_FIFO_blk[0] | proc_1_TLF_FIFO_blk[0] | proc_1_input_sync_blk[0] | proc_1_output_sync_blk[0]);
    assign proc_1_data_FIFO_blk[1] = 1'b0;
    assign proc_1_data_PIPO_blk[1] = 1'b0;
    assign proc_1_start_FIFO_blk[1] = 1'b0;
    assign proc_1_TLF_FIFO_blk[1] = 1'b0;
    assign proc_1_input_sync_blk[1] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_1_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_1[1] = dl_detect_out ? proc_dep_vld_vec_1_reg[1] : (proc_1_data_FIFO_blk[1] | proc_1_data_PIPO_blk[1] | proc_1_start_FIFO_blk[1] | proc_1_TLF_FIFO_blk[1] | proc_1_input_sync_blk[1] | proc_1_output_sync_blk[1]);
    assign proc_1_data_FIFO_blk[2] = 1'b0;
    assign proc_1_data_PIPO_blk[2] = 1'b0;
    assign proc_1_start_FIFO_blk[2] = 1'b0;
    assign proc_1_TLF_FIFO_blk[2] = 1'b0;
    assign proc_1_input_sync_blk[2] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_1_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_1[2] = dl_detect_out ? proc_dep_vld_vec_1_reg[2] : (proc_1_data_FIFO_blk[2] | proc_1_data_PIPO_blk[2] | proc_1_start_FIFO_blk[2] | proc_1_TLF_FIFO_blk[2] | proc_1_input_sync_blk[2] | proc_1_output_sync_blk[2]);
    assign proc_1_data_FIFO_blk[3] = 1'b0;
    assign proc_1_data_PIPO_blk[3] = 1'b0;
    assign proc_1_start_FIFO_blk[3] = 1'b0;
    assign proc_1_TLF_FIFO_blk[3] = 1'b0;
    assign proc_1_input_sync_blk[3] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_1_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_1[3] = dl_detect_out ? proc_dep_vld_vec_1_reg[3] : (proc_1_data_FIFO_blk[3] | proc_1_data_PIPO_blk[3] | proc_1_start_FIFO_blk[3] | proc_1_TLF_FIFO_blk[3] | proc_1_input_sync_blk[3] | proc_1_output_sync_blk[3]);
    assign proc_1_data_FIFO_blk[4] = 1'b0;
    assign proc_1_data_PIPO_blk[4] = 1'b0;
    assign proc_1_start_FIFO_blk[4] = 1'b0;
    assign proc_1_TLF_FIFO_blk[4] = 1'b0;
    assign proc_1_input_sync_blk[4] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_1_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_1[4] = dl_detect_out ? proc_dep_vld_vec_1_reg[4] : (proc_1_data_FIFO_blk[4] | proc_1_data_PIPO_blk[4] | proc_1_start_FIFO_blk[4] | proc_1_TLF_FIFO_blk[4] | proc_1_input_sync_blk[4] | proc_1_output_sync_blk[4]);
    assign proc_1_data_FIFO_blk[5] = 1'b0;
    assign proc_1_data_PIPO_blk[5] = 1'b0;
    assign proc_1_start_FIFO_blk[5] = 1'b0;
    assign proc_1_TLF_FIFO_blk[5] = 1'b0;
    assign proc_1_input_sync_blk[5] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_1_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_1[5] = dl_detect_out ? proc_dep_vld_vec_1_reg[5] : (proc_1_data_FIFO_blk[5] | proc_1_data_PIPO_blk[5] | proc_1_start_FIFO_blk[5] | proc_1_TLF_FIFO_blk[5] | proc_1_input_sync_blk[5] | proc_1_output_sync_blk[5]);
    assign proc_1_data_FIFO_blk[6] = 1'b0;
    assign proc_1_data_PIPO_blk[6] = 1'b0;
    assign proc_1_start_FIFO_blk[6] = 1'b0;
    assign proc_1_TLF_FIFO_blk[6] = 1'b0;
    assign proc_1_input_sync_blk[6] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_1_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_1[6] = dl_detect_out ? proc_dep_vld_vec_1_reg[6] : (proc_1_data_FIFO_blk[6] | proc_1_data_PIPO_blk[6] | proc_1_start_FIFO_blk[6] | proc_1_TLF_FIFO_blk[6] | proc_1_input_sync_blk[6] | proc_1_output_sync_blk[6]);
    assign proc_1_data_FIFO_blk[7] = 1'b0;
    assign proc_1_data_PIPO_blk[7] = 1'b0;
    assign proc_1_start_FIFO_blk[7] = 1'b0;
    assign proc_1_TLF_FIFO_blk[7] = 1'b0;
    assign proc_1_input_sync_blk[7] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_1_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_1[7] = dl_detect_out ? proc_dep_vld_vec_1_reg[7] : (proc_1_data_FIFO_blk[7] | proc_1_data_PIPO_blk[7] | proc_1_start_FIFO_blk[7] | proc_1_TLF_FIFO_blk[7] | proc_1_input_sync_blk[7] | proc_1_output_sync_blk[7]);
    assign proc_1_data_FIFO_blk[8] = 1'b0;
    assign proc_1_data_PIPO_blk[8] = 1'b0;
    assign proc_1_start_FIFO_blk[8] = 1'b0;
    assign proc_1_TLF_FIFO_blk[8] = 1'b0;
    assign proc_1_input_sync_blk[8] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_1_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_1[8] = dl_detect_out ? proc_dep_vld_vec_1_reg[8] : (proc_1_data_FIFO_blk[8] | proc_1_data_PIPO_blk[8] | proc_1_start_FIFO_blk[8] | proc_1_TLF_FIFO_blk[8] | proc_1_input_sync_blk[8] | proc_1_output_sync_blk[8]);
    assign proc_1_data_FIFO_blk[9] = 1'b0;
    assign proc_1_data_PIPO_blk[9] = 1'b0;
    assign proc_1_start_FIFO_blk[9] = 1'b0;
    assign proc_1_TLF_FIFO_blk[9] = 1'b0;
    assign proc_1_input_sync_blk[9] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_1_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_1[9] = dl_detect_out ? proc_dep_vld_vec_1_reg[9] : (proc_1_data_FIFO_blk[9] | proc_1_data_PIPO_blk[9] | proc_1_start_FIFO_blk[9] | proc_1_TLF_FIFO_blk[9] | proc_1_input_sync_blk[9] | proc_1_output_sync_blk[9]);
    assign proc_1_data_FIFO_blk[10] = 1'b0;
    assign proc_1_data_PIPO_blk[10] = 1'b0;
    assign proc_1_start_FIFO_blk[10] = 1'b0;
    assign proc_1_TLF_FIFO_blk[10] = 1'b0;
    assign proc_1_input_sync_blk[10] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_1_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_1[10] = dl_detect_out ? proc_dep_vld_vec_1_reg[10] : (proc_1_data_FIFO_blk[10] | proc_1_data_PIPO_blk[10] | proc_1_start_FIFO_blk[10] | proc_1_TLF_FIFO_blk[10] | proc_1_input_sync_blk[10] | proc_1_output_sync_blk[10]);
    assign proc_1_data_FIFO_blk[11] = 1'b0;
    assign proc_1_data_PIPO_blk[11] = 1'b0;
    assign proc_1_start_FIFO_blk[11] = 1'b0;
    assign proc_1_TLF_FIFO_blk[11] = 1'b0;
    assign proc_1_input_sync_blk[11] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_1_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_1[11] = dl_detect_out ? proc_dep_vld_vec_1_reg[11] : (proc_1_data_FIFO_blk[11] | proc_1_data_PIPO_blk[11] | proc_1_start_FIFO_blk[11] | proc_1_TLF_FIFO_blk[11] | proc_1_input_sync_blk[11] | proc_1_output_sync_blk[11]);
    assign proc_1_data_FIFO_blk[12] = 1'b0;
    assign proc_1_data_PIPO_blk[12] = 1'b0;
    assign proc_1_start_FIFO_blk[12] = 1'b0;
    assign proc_1_TLF_FIFO_blk[12] = 1'b0;
    assign proc_1_input_sync_blk[12] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_1_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_1[12] = dl_detect_out ? proc_dep_vld_vec_1_reg[12] : (proc_1_data_FIFO_blk[12] | proc_1_data_PIPO_blk[12] | proc_1_start_FIFO_blk[12] | proc_1_TLF_FIFO_blk[12] | proc_1_input_sync_blk[12] | proc_1_output_sync_blk[12]);
    assign proc_1_data_FIFO_blk[13] = 1'b0;
    assign proc_1_data_PIPO_blk[13] = 1'b0;
    assign proc_1_start_FIFO_blk[13] = 1'b0;
    assign proc_1_TLF_FIFO_blk[13] = 1'b0;
    assign proc_1_input_sync_blk[13] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_1_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_1[13] = dl_detect_out ? proc_dep_vld_vec_1_reg[13] : (proc_1_data_FIFO_blk[13] | proc_1_data_PIPO_blk[13] | proc_1_start_FIFO_blk[13] | proc_1_TLF_FIFO_blk[13] | proc_1_input_sync_blk[13] | proc_1_output_sync_blk[13]);
    assign proc_1_data_FIFO_blk[14] = 1'b0;
    assign proc_1_data_PIPO_blk[14] = 1'b0;
    assign proc_1_start_FIFO_blk[14] = 1'b0;
    assign proc_1_TLF_FIFO_blk[14] = 1'b0;
    assign proc_1_input_sync_blk[14] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_1_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_1[14] = dl_detect_out ? proc_dep_vld_vec_1_reg[14] : (proc_1_data_FIFO_blk[14] | proc_1_data_PIPO_blk[14] | proc_1_start_FIFO_blk[14] | proc_1_TLF_FIFO_blk[14] | proc_1_input_sync_blk[14] | proc_1_output_sync_blk[14]);
    assign proc_1_data_FIFO_blk[15] = 1'b0;
    assign proc_1_data_PIPO_blk[15] = 1'b0;
    assign proc_1_start_FIFO_blk[15] = 1'b0;
    assign proc_1_TLF_FIFO_blk[15] = 1'b0;
    assign proc_1_input_sync_blk[15] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_1_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_1[15] = dl_detect_out ? proc_dep_vld_vec_1_reg[15] : (proc_1_data_FIFO_blk[15] | proc_1_data_PIPO_blk[15] | proc_1_start_FIFO_blk[15] | proc_1_TLF_FIFO_blk[15] | proc_1_input_sync_blk[15] | proc_1_output_sync_blk[15]);
    assign proc_1_data_FIFO_blk[16] = 1'b0;
    assign proc_1_data_PIPO_blk[16] = 1'b0;
    assign proc_1_start_FIFO_blk[16] = 1'b0;
    assign proc_1_TLF_FIFO_blk[16] = 1'b0;
    assign proc_1_input_sync_blk[16] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_1_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_1[16] = dl_detect_out ? proc_dep_vld_vec_1_reg[16] : (proc_1_data_FIFO_blk[16] | proc_1_data_PIPO_blk[16] | proc_1_start_FIFO_blk[16] | proc_1_TLF_FIFO_blk[16] | proc_1_input_sync_blk[16] | proc_1_output_sync_blk[16]);
    assign proc_1_data_FIFO_blk[17] = 1'b0;
    assign proc_1_data_PIPO_blk[17] = 1'b0;
    assign proc_1_start_FIFO_blk[17] = 1'b0;
    assign proc_1_TLF_FIFO_blk[17] = 1'b0;
    assign proc_1_input_sync_blk[17] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_1_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_1[17] = dl_detect_out ? proc_dep_vld_vec_1_reg[17] : (proc_1_data_FIFO_blk[17] | proc_1_data_PIPO_blk[17] | proc_1_start_FIFO_blk[17] | proc_1_TLF_FIFO_blk[17] | proc_1_input_sync_blk[17] | proc_1_output_sync_blk[17]);
    assign proc_1_data_FIFO_blk[18] = 1'b0;
    assign proc_1_data_PIPO_blk[18] = 1'b0;
    assign proc_1_start_FIFO_blk[18] = 1'b0;
    assign proc_1_TLF_FIFO_blk[18] = 1'b0;
    assign proc_1_input_sync_blk[18] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_1_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_1[18] = dl_detect_out ? proc_dep_vld_vec_1_reg[18] : (proc_1_data_FIFO_blk[18] | proc_1_data_PIPO_blk[18] | proc_1_start_FIFO_blk[18] | proc_1_TLF_FIFO_blk[18] | proc_1_input_sync_blk[18] | proc_1_output_sync_blk[18]);
    assign proc_1_data_FIFO_blk[19] = 1'b0;
    assign proc_1_data_PIPO_blk[19] = 1'b0;
    assign proc_1_start_FIFO_blk[19] = 1'b0;
    assign proc_1_TLF_FIFO_blk[19] = 1'b0;
    assign proc_1_input_sync_blk[19] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_1_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_1[19] = dl_detect_out ? proc_dep_vld_vec_1_reg[19] : (proc_1_data_FIFO_blk[19] | proc_1_data_PIPO_blk[19] | proc_1_start_FIFO_blk[19] | proc_1_TLF_FIFO_blk[19] | proc_1_input_sync_blk[19] | proc_1_output_sync_blk[19]);
    assign proc_1_data_FIFO_blk[20] = 1'b0;
    assign proc_1_data_PIPO_blk[20] = 1'b0;
    assign proc_1_start_FIFO_blk[20] = 1'b0;
    assign proc_1_TLF_FIFO_blk[20] = 1'b0;
    assign proc_1_input_sync_blk[20] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_1_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_1[20] = dl_detect_out ? proc_dep_vld_vec_1_reg[20] : (proc_1_data_FIFO_blk[20] | proc_1_data_PIPO_blk[20] | proc_1_start_FIFO_blk[20] | proc_1_TLF_FIFO_blk[20] | proc_1_input_sync_blk[20] | proc_1_output_sync_blk[20]);
    assign proc_1_data_FIFO_blk[21] = 1'b0;
    assign proc_1_data_PIPO_blk[21] = 1'b0;
    assign proc_1_start_FIFO_blk[21] = 1'b0;
    assign proc_1_TLF_FIFO_blk[21] = 1'b0;
    assign proc_1_input_sync_blk[21] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_1_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_1[21] = dl_detect_out ? proc_dep_vld_vec_1_reg[21] : (proc_1_data_FIFO_blk[21] | proc_1_data_PIPO_blk[21] | proc_1_start_FIFO_blk[21] | proc_1_TLF_FIFO_blk[21] | proc_1_input_sync_blk[21] | proc_1_output_sync_blk[21]);
    assign proc_1_data_FIFO_blk[22] = 1'b0;
    assign proc_1_data_PIPO_blk[22] = 1'b0;
    assign proc_1_start_FIFO_blk[22] = 1'b0;
    assign proc_1_TLF_FIFO_blk[22] = 1'b0;
    assign proc_1_input_sync_blk[22] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_1_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_1[22] = dl_detect_out ? proc_dep_vld_vec_1_reg[22] : (proc_1_data_FIFO_blk[22] | proc_1_data_PIPO_blk[22] | proc_1_start_FIFO_blk[22] | proc_1_TLF_FIFO_blk[22] | proc_1_input_sync_blk[22] | proc_1_output_sync_blk[22]);
    assign proc_1_data_FIFO_blk[23] = 1'b0;
    assign proc_1_data_PIPO_blk[23] = 1'b0;
    assign proc_1_start_FIFO_blk[23] = 1'b0;
    assign proc_1_TLF_FIFO_blk[23] = 1'b0;
    assign proc_1_input_sync_blk[23] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_1_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_1[23] = dl_detect_out ? proc_dep_vld_vec_1_reg[23] : (proc_1_data_FIFO_blk[23] | proc_1_data_PIPO_blk[23] | proc_1_start_FIFO_blk[23] | proc_1_TLF_FIFO_blk[23] | proc_1_input_sync_blk[23] | proc_1_output_sync_blk[23]);
    assign proc_1_data_FIFO_blk[24] = 1'b0;
    assign proc_1_data_PIPO_blk[24] = 1'b0;
    assign proc_1_start_FIFO_blk[24] = 1'b0;
    assign proc_1_TLF_FIFO_blk[24] = 1'b0;
    assign proc_1_input_sync_blk[24] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_1_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_1[24] = dl_detect_out ? proc_dep_vld_vec_1_reg[24] : (proc_1_data_FIFO_blk[24] | proc_1_data_PIPO_blk[24] | proc_1_start_FIFO_blk[24] | proc_1_TLF_FIFO_blk[24] | proc_1_input_sync_blk[24] | proc_1_output_sync_blk[24]);
    assign proc_1_data_FIFO_blk[25] = 1'b0;
    assign proc_1_data_PIPO_blk[25] = 1'b0;
    assign proc_1_start_FIFO_blk[25] = 1'b0;
    assign proc_1_TLF_FIFO_blk[25] = 1'b0;
    assign proc_1_input_sync_blk[25] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_1_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_1[25] = dl_detect_out ? proc_dep_vld_vec_1_reg[25] : (proc_1_data_FIFO_blk[25] | proc_1_data_PIPO_blk[25] | proc_1_start_FIFO_blk[25] | proc_1_TLF_FIFO_blk[25] | proc_1_input_sync_blk[25] | proc_1_output_sync_blk[25]);
    assign proc_1_data_FIFO_blk[26] = 1'b0;
    assign proc_1_data_PIPO_blk[26] = 1'b0;
    assign proc_1_start_FIFO_blk[26] = 1'b0;
    assign proc_1_TLF_FIFO_blk[26] = 1'b0;
    assign proc_1_input_sync_blk[26] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_1_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_1[26] = dl_detect_out ? proc_dep_vld_vec_1_reg[26] : (proc_1_data_FIFO_blk[26] | proc_1_data_PIPO_blk[26] | proc_1_start_FIFO_blk[26] | proc_1_TLF_FIFO_blk[26] | proc_1_input_sync_blk[26] | proc_1_output_sync_blk[26]);
    assign proc_1_data_FIFO_blk[27] = 1'b0;
    assign proc_1_data_PIPO_blk[27] = 1'b0;
    assign proc_1_start_FIFO_blk[27] = 1'b0;
    assign proc_1_TLF_FIFO_blk[27] = 1'b0;
    assign proc_1_input_sync_blk[27] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_1_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_1[27] = dl_detect_out ? proc_dep_vld_vec_1_reg[27] : (proc_1_data_FIFO_blk[27] | proc_1_data_PIPO_blk[27] | proc_1_start_FIFO_blk[27] | proc_1_TLF_FIFO_blk[27] | proc_1_input_sync_blk[27] | proc_1_output_sync_blk[27]);
    assign proc_1_data_FIFO_blk[28] = 1'b0;
    assign proc_1_data_PIPO_blk[28] = 1'b0;
    assign proc_1_start_FIFO_blk[28] = 1'b0;
    assign proc_1_TLF_FIFO_blk[28] = 1'b0;
    assign proc_1_input_sync_blk[28] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_1_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_1[28] = dl_detect_out ? proc_dep_vld_vec_1_reg[28] : (proc_1_data_FIFO_blk[28] | proc_1_data_PIPO_blk[28] | proc_1_start_FIFO_blk[28] | proc_1_TLF_FIFO_blk[28] | proc_1_input_sync_blk[28] | proc_1_output_sync_blk[28]);
    assign proc_1_data_FIFO_blk[29] = 1'b0;
    assign proc_1_data_PIPO_blk[29] = 1'b0;
    assign proc_1_start_FIFO_blk[29] = 1'b0;
    assign proc_1_TLF_FIFO_blk[29] = 1'b0;
    assign proc_1_input_sync_blk[29] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_1_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_1[29] = dl_detect_out ? proc_dep_vld_vec_1_reg[29] : (proc_1_data_FIFO_blk[29] | proc_1_data_PIPO_blk[29] | proc_1_start_FIFO_blk[29] | proc_1_TLF_FIFO_blk[29] | proc_1_input_sync_blk[29] | proc_1_output_sync_blk[29]);
    assign proc_1_data_FIFO_blk[30] = 1'b0;
    assign proc_1_data_PIPO_blk[30] = 1'b0;
    assign proc_1_start_FIFO_blk[30] = 1'b0;
    assign proc_1_TLF_FIFO_blk[30] = 1'b0;
    assign proc_1_input_sync_blk[30] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_1_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_1[30] = dl_detect_out ? proc_dep_vld_vec_1_reg[30] : (proc_1_data_FIFO_blk[30] | proc_1_data_PIPO_blk[30] | proc_1_start_FIFO_blk[30] | proc_1_TLF_FIFO_blk[30] | proc_1_input_sync_blk[30] | proc_1_output_sync_blk[30]);
    assign proc_1_data_FIFO_blk[31] = 1'b0;
    assign proc_1_data_PIPO_blk[31] = 1'b0;
    assign proc_1_start_FIFO_blk[31] = 1'b0;
    assign proc_1_TLF_FIFO_blk[31] = 1'b0;
    assign proc_1_input_sync_blk[31] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_1_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_1[31] = dl_detect_out ? proc_dep_vld_vec_1_reg[31] : (proc_1_data_FIFO_blk[31] | proc_1_data_PIPO_blk[31] | proc_1_start_FIFO_blk[31] | proc_1_TLF_FIFO_blk[31] | proc_1_input_sync_blk[31] | proc_1_output_sync_blk[31]);
    assign proc_1_data_FIFO_blk[32] = 1'b0;
    assign proc_1_data_PIPO_blk[32] = 1'b0;
    assign proc_1_start_FIFO_blk[32] = 1'b0;
    assign proc_1_TLF_FIFO_blk[32] = 1'b0;
    assign proc_1_input_sync_blk[32] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_1_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_1[32] = dl_detect_out ? proc_dep_vld_vec_1_reg[32] : (proc_1_data_FIFO_blk[32] | proc_1_data_PIPO_blk[32] | proc_1_start_FIFO_blk[32] | proc_1_TLF_FIFO_blk[32] | proc_1_input_sync_blk[32] | proc_1_output_sync_blk[32]);
    assign proc_1_data_FIFO_blk[33] = 1'b0;
    assign proc_1_data_PIPO_blk[33] = 1'b0;
    assign proc_1_start_FIFO_blk[33] = 1'b0;
    assign proc_1_TLF_FIFO_blk[33] = 1'b0;
    assign proc_1_input_sync_blk[33] = 1'b0 | (ap_sync_ReadA_U0_ap_ready & ReadA_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_1_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_1[33] = dl_detect_out ? proc_dep_vld_vec_1_reg[33] : (proc_1_data_FIFO_blk[33] | proc_1_data_PIPO_blk[33] | proc_1_start_FIFO_blk[33] | proc_1_TLF_FIFO_blk[33] | proc_1_input_sync_blk[33] | proc_1_output_sync_blk[33]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_1_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_1_reg <= proc_dep_vld_vec_1;
        end
    end
    assign in_chan_dep_vld_vec_1[0] = dep_chan_vld_0_1;
    assign in_chan_dep_data_vec_1[39 : 0] = dep_chan_data_0_1;
    assign token_in_vec_1[0] = token_0_1;
    assign in_chan_dep_vld_vec_1[1] = dep_chan_vld_2_1;
    assign in_chan_dep_data_vec_1[79 : 40] = dep_chan_data_2_1;
    assign token_in_vec_1[1] = token_2_1;
    assign in_chan_dep_vld_vec_1[2] = dep_chan_vld_3_1;
    assign in_chan_dep_data_vec_1[119 : 80] = dep_chan_data_3_1;
    assign token_in_vec_1[2] = token_3_1;
    assign in_chan_dep_vld_vec_1[3] = dep_chan_vld_6_1;
    assign in_chan_dep_data_vec_1[159 : 120] = dep_chan_data_6_1;
    assign token_in_vec_1[3] = token_6_1;
    assign in_chan_dep_vld_vec_1[4] = dep_chan_vld_7_1;
    assign in_chan_dep_data_vec_1[199 : 160] = dep_chan_data_7_1;
    assign token_in_vec_1[4] = token_7_1;
    assign in_chan_dep_vld_vec_1[5] = dep_chan_vld_8_1;
    assign in_chan_dep_data_vec_1[239 : 200] = dep_chan_data_8_1;
    assign token_in_vec_1[5] = token_8_1;
    assign in_chan_dep_vld_vec_1[6] = dep_chan_vld_9_1;
    assign in_chan_dep_data_vec_1[279 : 240] = dep_chan_data_9_1;
    assign token_in_vec_1[6] = token_9_1;
    assign in_chan_dep_vld_vec_1[7] = dep_chan_vld_10_1;
    assign in_chan_dep_data_vec_1[319 : 280] = dep_chan_data_10_1;
    assign token_in_vec_1[7] = token_10_1;
    assign in_chan_dep_vld_vec_1[8] = dep_chan_vld_11_1;
    assign in_chan_dep_data_vec_1[359 : 320] = dep_chan_data_11_1;
    assign token_in_vec_1[8] = token_11_1;
    assign in_chan_dep_vld_vec_1[9] = dep_chan_vld_12_1;
    assign in_chan_dep_data_vec_1[399 : 360] = dep_chan_data_12_1;
    assign token_in_vec_1[9] = token_12_1;
    assign in_chan_dep_vld_vec_1[10] = dep_chan_vld_13_1;
    assign in_chan_dep_data_vec_1[439 : 400] = dep_chan_data_13_1;
    assign token_in_vec_1[10] = token_13_1;
    assign in_chan_dep_vld_vec_1[11] = dep_chan_vld_14_1;
    assign in_chan_dep_data_vec_1[479 : 440] = dep_chan_data_14_1;
    assign token_in_vec_1[11] = token_14_1;
    assign in_chan_dep_vld_vec_1[12] = dep_chan_vld_15_1;
    assign in_chan_dep_data_vec_1[519 : 480] = dep_chan_data_15_1;
    assign token_in_vec_1[12] = token_15_1;
    assign in_chan_dep_vld_vec_1[13] = dep_chan_vld_16_1;
    assign in_chan_dep_data_vec_1[559 : 520] = dep_chan_data_16_1;
    assign token_in_vec_1[13] = token_16_1;
    assign in_chan_dep_vld_vec_1[14] = dep_chan_vld_17_1;
    assign in_chan_dep_data_vec_1[599 : 560] = dep_chan_data_17_1;
    assign token_in_vec_1[14] = token_17_1;
    assign in_chan_dep_vld_vec_1[15] = dep_chan_vld_18_1;
    assign in_chan_dep_data_vec_1[639 : 600] = dep_chan_data_18_1;
    assign token_in_vec_1[15] = token_18_1;
    assign in_chan_dep_vld_vec_1[16] = dep_chan_vld_19_1;
    assign in_chan_dep_data_vec_1[679 : 640] = dep_chan_data_19_1;
    assign token_in_vec_1[16] = token_19_1;
    assign in_chan_dep_vld_vec_1[17] = dep_chan_vld_20_1;
    assign in_chan_dep_data_vec_1[719 : 680] = dep_chan_data_20_1;
    assign token_in_vec_1[17] = token_20_1;
    assign in_chan_dep_vld_vec_1[18] = dep_chan_vld_21_1;
    assign in_chan_dep_data_vec_1[759 : 720] = dep_chan_data_21_1;
    assign token_in_vec_1[18] = token_21_1;
    assign in_chan_dep_vld_vec_1[19] = dep_chan_vld_22_1;
    assign in_chan_dep_data_vec_1[799 : 760] = dep_chan_data_22_1;
    assign token_in_vec_1[19] = token_22_1;
    assign in_chan_dep_vld_vec_1[20] = dep_chan_vld_23_1;
    assign in_chan_dep_data_vec_1[839 : 800] = dep_chan_data_23_1;
    assign token_in_vec_1[20] = token_23_1;
    assign in_chan_dep_vld_vec_1[21] = dep_chan_vld_24_1;
    assign in_chan_dep_data_vec_1[879 : 840] = dep_chan_data_24_1;
    assign token_in_vec_1[21] = token_24_1;
    assign in_chan_dep_vld_vec_1[22] = dep_chan_vld_25_1;
    assign in_chan_dep_data_vec_1[919 : 880] = dep_chan_data_25_1;
    assign token_in_vec_1[22] = token_25_1;
    assign in_chan_dep_vld_vec_1[23] = dep_chan_vld_26_1;
    assign in_chan_dep_data_vec_1[959 : 920] = dep_chan_data_26_1;
    assign token_in_vec_1[23] = token_26_1;
    assign in_chan_dep_vld_vec_1[24] = dep_chan_vld_27_1;
    assign in_chan_dep_data_vec_1[999 : 960] = dep_chan_data_27_1;
    assign token_in_vec_1[24] = token_27_1;
    assign in_chan_dep_vld_vec_1[25] = dep_chan_vld_28_1;
    assign in_chan_dep_data_vec_1[1039 : 1000] = dep_chan_data_28_1;
    assign token_in_vec_1[25] = token_28_1;
    assign in_chan_dep_vld_vec_1[26] = dep_chan_vld_29_1;
    assign in_chan_dep_data_vec_1[1079 : 1040] = dep_chan_data_29_1;
    assign token_in_vec_1[26] = token_29_1;
    assign in_chan_dep_vld_vec_1[27] = dep_chan_vld_30_1;
    assign in_chan_dep_data_vec_1[1119 : 1080] = dep_chan_data_30_1;
    assign token_in_vec_1[27] = token_30_1;
    assign in_chan_dep_vld_vec_1[28] = dep_chan_vld_31_1;
    assign in_chan_dep_data_vec_1[1159 : 1120] = dep_chan_data_31_1;
    assign token_in_vec_1[28] = token_31_1;
    assign in_chan_dep_vld_vec_1[29] = dep_chan_vld_32_1;
    assign in_chan_dep_data_vec_1[1199 : 1160] = dep_chan_data_32_1;
    assign token_in_vec_1[29] = token_32_1;
    assign in_chan_dep_vld_vec_1[30] = dep_chan_vld_33_1;
    assign in_chan_dep_data_vec_1[1239 : 1200] = dep_chan_data_33_1;
    assign token_in_vec_1[30] = token_33_1;
    assign in_chan_dep_vld_vec_1[31] = dep_chan_vld_34_1;
    assign in_chan_dep_data_vec_1[1279 : 1240] = dep_chan_data_34_1;
    assign token_in_vec_1[31] = token_34_1;
    assign in_chan_dep_vld_vec_1[32] = dep_chan_vld_35_1;
    assign in_chan_dep_data_vec_1[1319 : 1280] = dep_chan_data_35_1;
    assign token_in_vec_1[32] = token_35_1;
    assign in_chan_dep_vld_vec_1[33] = dep_chan_vld_36_1;
    assign in_chan_dep_data_vec_1[1359 : 1320] = dep_chan_data_36_1;
    assign token_in_vec_1[33] = token_36_1;
    assign dep_chan_vld_1_2 = out_chan_dep_vld_vec_1[0];
    assign dep_chan_data_1_2 = out_chan_dep_data_1;
    assign token_1_2 = token_out_vec_1[0];
    assign dep_chan_vld_1_0 = out_chan_dep_vld_vec_1[1];
    assign dep_chan_data_1_0 = out_chan_dep_data_1;
    assign token_1_0 = token_out_vec_1[1];
    assign dep_chan_vld_1_3 = out_chan_dep_vld_vec_1[2];
    assign dep_chan_data_1_3 = out_chan_dep_data_1;
    assign token_1_3 = token_out_vec_1[2];
    assign dep_chan_vld_1_6 = out_chan_dep_vld_vec_1[3];
    assign dep_chan_data_1_6 = out_chan_dep_data_1;
    assign token_1_6 = token_out_vec_1[3];
    assign dep_chan_vld_1_7 = out_chan_dep_vld_vec_1[4];
    assign dep_chan_data_1_7 = out_chan_dep_data_1;
    assign token_1_7 = token_out_vec_1[4];
    assign dep_chan_vld_1_8 = out_chan_dep_vld_vec_1[5];
    assign dep_chan_data_1_8 = out_chan_dep_data_1;
    assign token_1_8 = token_out_vec_1[5];
    assign dep_chan_vld_1_9 = out_chan_dep_vld_vec_1[6];
    assign dep_chan_data_1_9 = out_chan_dep_data_1;
    assign token_1_9 = token_out_vec_1[6];
    assign dep_chan_vld_1_10 = out_chan_dep_vld_vec_1[7];
    assign dep_chan_data_1_10 = out_chan_dep_data_1;
    assign token_1_10 = token_out_vec_1[7];
    assign dep_chan_vld_1_11 = out_chan_dep_vld_vec_1[8];
    assign dep_chan_data_1_11 = out_chan_dep_data_1;
    assign token_1_11 = token_out_vec_1[8];
    assign dep_chan_vld_1_12 = out_chan_dep_vld_vec_1[9];
    assign dep_chan_data_1_12 = out_chan_dep_data_1;
    assign token_1_12 = token_out_vec_1[9];
    assign dep_chan_vld_1_13 = out_chan_dep_vld_vec_1[10];
    assign dep_chan_data_1_13 = out_chan_dep_data_1;
    assign token_1_13 = token_out_vec_1[10];
    assign dep_chan_vld_1_14 = out_chan_dep_vld_vec_1[11];
    assign dep_chan_data_1_14 = out_chan_dep_data_1;
    assign token_1_14 = token_out_vec_1[11];
    assign dep_chan_vld_1_15 = out_chan_dep_vld_vec_1[12];
    assign dep_chan_data_1_15 = out_chan_dep_data_1;
    assign token_1_15 = token_out_vec_1[12];
    assign dep_chan_vld_1_16 = out_chan_dep_vld_vec_1[13];
    assign dep_chan_data_1_16 = out_chan_dep_data_1;
    assign token_1_16 = token_out_vec_1[13];
    assign dep_chan_vld_1_17 = out_chan_dep_vld_vec_1[14];
    assign dep_chan_data_1_17 = out_chan_dep_data_1;
    assign token_1_17 = token_out_vec_1[14];
    assign dep_chan_vld_1_18 = out_chan_dep_vld_vec_1[15];
    assign dep_chan_data_1_18 = out_chan_dep_data_1;
    assign token_1_18 = token_out_vec_1[15];
    assign dep_chan_vld_1_19 = out_chan_dep_vld_vec_1[16];
    assign dep_chan_data_1_19 = out_chan_dep_data_1;
    assign token_1_19 = token_out_vec_1[16];
    assign dep_chan_vld_1_20 = out_chan_dep_vld_vec_1[17];
    assign dep_chan_data_1_20 = out_chan_dep_data_1;
    assign token_1_20 = token_out_vec_1[17];
    assign dep_chan_vld_1_21 = out_chan_dep_vld_vec_1[18];
    assign dep_chan_data_1_21 = out_chan_dep_data_1;
    assign token_1_21 = token_out_vec_1[18];
    assign dep_chan_vld_1_22 = out_chan_dep_vld_vec_1[19];
    assign dep_chan_data_1_22 = out_chan_dep_data_1;
    assign token_1_22 = token_out_vec_1[19];
    assign dep_chan_vld_1_23 = out_chan_dep_vld_vec_1[20];
    assign dep_chan_data_1_23 = out_chan_dep_data_1;
    assign token_1_23 = token_out_vec_1[20];
    assign dep_chan_vld_1_24 = out_chan_dep_vld_vec_1[21];
    assign dep_chan_data_1_24 = out_chan_dep_data_1;
    assign token_1_24 = token_out_vec_1[21];
    assign dep_chan_vld_1_25 = out_chan_dep_vld_vec_1[22];
    assign dep_chan_data_1_25 = out_chan_dep_data_1;
    assign token_1_25 = token_out_vec_1[22];
    assign dep_chan_vld_1_26 = out_chan_dep_vld_vec_1[23];
    assign dep_chan_data_1_26 = out_chan_dep_data_1;
    assign token_1_26 = token_out_vec_1[23];
    assign dep_chan_vld_1_27 = out_chan_dep_vld_vec_1[24];
    assign dep_chan_data_1_27 = out_chan_dep_data_1;
    assign token_1_27 = token_out_vec_1[24];
    assign dep_chan_vld_1_28 = out_chan_dep_vld_vec_1[25];
    assign dep_chan_data_1_28 = out_chan_dep_data_1;
    assign token_1_28 = token_out_vec_1[25];
    assign dep_chan_vld_1_29 = out_chan_dep_vld_vec_1[26];
    assign dep_chan_data_1_29 = out_chan_dep_data_1;
    assign token_1_29 = token_out_vec_1[26];
    assign dep_chan_vld_1_30 = out_chan_dep_vld_vec_1[27];
    assign dep_chan_data_1_30 = out_chan_dep_data_1;
    assign token_1_30 = token_out_vec_1[27];
    assign dep_chan_vld_1_31 = out_chan_dep_vld_vec_1[28];
    assign dep_chan_data_1_31 = out_chan_dep_data_1;
    assign token_1_31 = token_out_vec_1[28];
    assign dep_chan_vld_1_32 = out_chan_dep_vld_vec_1[29];
    assign dep_chan_data_1_32 = out_chan_dep_data_1;
    assign token_1_32 = token_out_vec_1[29];
    assign dep_chan_vld_1_33 = out_chan_dep_vld_vec_1[30];
    assign dep_chan_data_1_33 = out_chan_dep_data_1;
    assign token_1_33 = token_out_vec_1[30];
    assign dep_chan_vld_1_34 = out_chan_dep_vld_vec_1[31];
    assign dep_chan_data_1_34 = out_chan_dep_data_1;
    assign token_1_34 = token_out_vec_1[31];
    assign dep_chan_vld_1_35 = out_chan_dep_vld_vec_1[32];
    assign dep_chan_data_1_35 = out_chan_dep_data_1;
    assign token_1_35 = token_out_vec_1[32];
    assign dep_chan_vld_1_36 = out_chan_dep_vld_vec_1[33];
    assign dep_chan_data_1_36 = out_chan_dep_data_1;
    assign token_1_36 = token_out_vec_1[33];

    // Process: TransposeA_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 2, 2, 2) MatrixMultiplicationKernel_hls_deadlock_detect_unit_2 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_2),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_2),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_2),
        .token_in_vec(token_in_vec_2),
        .dl_detect_in(dl_detect_out),
        .origin(origin[2]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_2),
        .out_chan_dep_data(out_chan_dep_data_2),
        .token_out_vec(token_out_vec_2),
        .dl_detect_out(dl_in_vec[2]));

    assign proc_2_data_FIFO_blk[0] = 1'b0 | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_0_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_1_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_2_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_3_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_4_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_5_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_6_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_7_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_8_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_9_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_10_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_11_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_12_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_13_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_14_blk_n) | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aSplit_15_blk_n) | (~TransposeA_U0.size_n_blk_n) | (~TransposeA_U0.size_k_blk_n) | (~TransposeA_U0.size_m_blk_n);
    assign proc_2_data_PIPO_blk[0] = 1'b0;
    assign proc_2_start_FIFO_blk[0] = 1'b0 | (~start_for_TransposeA_U0_U.if_empty_n & TransposeA_U0.ap_idle & ~start_for_TransposeA_U0_U.if_write);
    assign proc_2_TLF_FIFO_blk[0] = 1'b0;
    assign proc_2_input_sync_blk[0] = 1'b0;
    assign proc_2_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_2[0] = dl_detect_out ? proc_dep_vld_vec_2_reg[0] : (proc_2_data_FIFO_blk[0] | proc_2_data_PIPO_blk[0] | proc_2_start_FIFO_blk[0] | proc_2_TLF_FIFO_blk[0] | proc_2_input_sync_blk[0] | proc_2_output_sync_blk[0]);
    assign proc_2_data_FIFO_blk[1] = 1'b0 | (~TransposeA_U0.grp_TransposeA_Pipeline_TransposeA_N0_TransposeA_M0_TransposeA_K_VITIS_LOOP_153_1_fu_96.aPipes_0_blk_n);
    assign proc_2_data_PIPO_blk[1] = 1'b0;
    assign proc_2_start_FIFO_blk[1] = 1'b0;
    assign proc_2_TLF_FIFO_blk[1] = 1'b0;
    assign proc_2_input_sync_blk[1] = 1'b0;
    assign proc_2_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_2[1] = dl_detect_out ? proc_dep_vld_vec_2_reg[1] : (proc_2_data_FIFO_blk[1] | proc_2_data_PIPO_blk[1] | proc_2_start_FIFO_blk[1] | proc_2_TLF_FIFO_blk[1] | proc_2_input_sync_blk[1] | proc_2_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_2_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_2_reg <= proc_dep_vld_vec_2;
        end
    end
    assign in_chan_dep_vld_vec_2[0] = dep_chan_vld_1_2;
    assign in_chan_dep_data_vec_2[39 : 0] = dep_chan_data_1_2;
    assign token_in_vec_2[0] = token_1_2;
    assign in_chan_dep_vld_vec_2[1] = dep_chan_vld_6_2;
    assign in_chan_dep_data_vec_2[79 : 40] = dep_chan_data_6_2;
    assign token_in_vec_2[1] = token_6_2;
    assign dep_chan_vld_2_1 = out_chan_dep_vld_vec_2[0];
    assign dep_chan_data_2_1 = out_chan_dep_data_2;
    assign token_2_1 = token_out_vec_2[0];
    assign dep_chan_vld_2_6 = out_chan_dep_vld_vec_2[1];
    assign dep_chan_data_2_6 = out_chan_dep_data_2;
    assign token_2_6 = token_out_vec_2[1];

    // Process: ReadB_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 3, 34, 34) MatrixMultiplicationKernel_hls_deadlock_detect_unit_3 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_3),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_3),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_3),
        .token_in_vec(token_in_vec_3),
        .dl_detect_in(dl_detect_out),
        .origin(origin[3]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_3),
        .out_chan_dep_data(out_chan_dep_data_3),
        .token_out_vec(token_out_vec_3),
        .dl_detect_out(dl_in_vec[3]));

    assign proc_3_data_FIFO_blk[0] = 1'b0 | (~ReadB_U0.grp_ReadB_Pipeline_ReadB_OuterTile_N_ReadB_OuterTile_M_ReadB_K_ReadB_BufferB_M1_fu_122.bMemory_blk_n) | (~ReadB_U0.size_n_c4_blk_n) | (~ReadB_U0.size_k_c7_blk_n) | (~ReadB_U0.size_m_c12_blk_n);
    assign proc_3_data_PIPO_blk[0] = 1'b0;
    assign proc_3_start_FIFO_blk[0] = 1'b0 | (~start_for_ConvertWidthB_U0_U.if_full_n & ReadB_U0.ap_start & ~ReadB_U0.real_start & (trans_in_cnt_1 == trans_out_cnt_1) & ~start_for_ConvertWidthB_U0_U.if_read);
    assign proc_3_TLF_FIFO_blk[0] = 1'b0;
    assign proc_3_input_sync_blk[0] = 1'b0;
    assign proc_3_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_3[0] = dl_detect_out ? proc_dep_vld_vec_3_reg[0] : (proc_3_data_FIFO_blk[0] | proc_3_data_PIPO_blk[0] | proc_3_start_FIFO_blk[0] | proc_3_TLF_FIFO_blk[0] | proc_3_input_sync_blk[0] | proc_3_output_sync_blk[0]);
    assign proc_3_data_FIFO_blk[1] = 1'b0;
    assign proc_3_data_PIPO_blk[1] = 1'b0;
    assign proc_3_start_FIFO_blk[1] = 1'b0;
    assign proc_3_TLF_FIFO_blk[1] = 1'b0;
    assign proc_3_input_sync_blk[1] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_3_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_3[1] = dl_detect_out ? proc_dep_vld_vec_3_reg[1] : (proc_3_data_FIFO_blk[1] | proc_3_data_PIPO_blk[1] | proc_3_start_FIFO_blk[1] | proc_3_TLF_FIFO_blk[1] | proc_3_input_sync_blk[1] | proc_3_output_sync_blk[1]);
    assign proc_3_data_FIFO_blk[2] = 1'b0;
    assign proc_3_data_PIPO_blk[2] = 1'b0;
    assign proc_3_start_FIFO_blk[2] = 1'b0;
    assign proc_3_TLF_FIFO_blk[2] = 1'b0;
    assign proc_3_input_sync_blk[2] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_3_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_3[2] = dl_detect_out ? proc_dep_vld_vec_3_reg[2] : (proc_3_data_FIFO_blk[2] | proc_3_data_PIPO_blk[2] | proc_3_start_FIFO_blk[2] | proc_3_TLF_FIFO_blk[2] | proc_3_input_sync_blk[2] | proc_3_output_sync_blk[2]);
    assign proc_3_data_FIFO_blk[3] = 1'b0;
    assign proc_3_data_PIPO_blk[3] = 1'b0;
    assign proc_3_start_FIFO_blk[3] = 1'b0;
    assign proc_3_TLF_FIFO_blk[3] = 1'b0;
    assign proc_3_input_sync_blk[3] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_3_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_3[3] = dl_detect_out ? proc_dep_vld_vec_3_reg[3] : (proc_3_data_FIFO_blk[3] | proc_3_data_PIPO_blk[3] | proc_3_start_FIFO_blk[3] | proc_3_TLF_FIFO_blk[3] | proc_3_input_sync_blk[3] | proc_3_output_sync_blk[3]);
    assign proc_3_data_FIFO_blk[4] = 1'b0;
    assign proc_3_data_PIPO_blk[4] = 1'b0;
    assign proc_3_start_FIFO_blk[4] = 1'b0;
    assign proc_3_TLF_FIFO_blk[4] = 1'b0;
    assign proc_3_input_sync_blk[4] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_3_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_3[4] = dl_detect_out ? proc_dep_vld_vec_3_reg[4] : (proc_3_data_FIFO_blk[4] | proc_3_data_PIPO_blk[4] | proc_3_start_FIFO_blk[4] | proc_3_TLF_FIFO_blk[4] | proc_3_input_sync_blk[4] | proc_3_output_sync_blk[4]);
    assign proc_3_data_FIFO_blk[5] = 1'b0;
    assign proc_3_data_PIPO_blk[5] = 1'b0;
    assign proc_3_start_FIFO_blk[5] = 1'b0;
    assign proc_3_TLF_FIFO_blk[5] = 1'b0;
    assign proc_3_input_sync_blk[5] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_3_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_3[5] = dl_detect_out ? proc_dep_vld_vec_3_reg[5] : (proc_3_data_FIFO_blk[5] | proc_3_data_PIPO_blk[5] | proc_3_start_FIFO_blk[5] | proc_3_TLF_FIFO_blk[5] | proc_3_input_sync_blk[5] | proc_3_output_sync_blk[5]);
    assign proc_3_data_FIFO_blk[6] = 1'b0;
    assign proc_3_data_PIPO_blk[6] = 1'b0;
    assign proc_3_start_FIFO_blk[6] = 1'b0;
    assign proc_3_TLF_FIFO_blk[6] = 1'b0;
    assign proc_3_input_sync_blk[6] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_3_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_3[6] = dl_detect_out ? proc_dep_vld_vec_3_reg[6] : (proc_3_data_FIFO_blk[6] | proc_3_data_PIPO_blk[6] | proc_3_start_FIFO_blk[6] | proc_3_TLF_FIFO_blk[6] | proc_3_input_sync_blk[6] | proc_3_output_sync_blk[6]);
    assign proc_3_data_FIFO_blk[7] = 1'b0;
    assign proc_3_data_PIPO_blk[7] = 1'b0;
    assign proc_3_start_FIFO_blk[7] = 1'b0;
    assign proc_3_TLF_FIFO_blk[7] = 1'b0;
    assign proc_3_input_sync_blk[7] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_3_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_3[7] = dl_detect_out ? proc_dep_vld_vec_3_reg[7] : (proc_3_data_FIFO_blk[7] | proc_3_data_PIPO_blk[7] | proc_3_start_FIFO_blk[7] | proc_3_TLF_FIFO_blk[7] | proc_3_input_sync_blk[7] | proc_3_output_sync_blk[7]);
    assign proc_3_data_FIFO_blk[8] = 1'b0;
    assign proc_3_data_PIPO_blk[8] = 1'b0;
    assign proc_3_start_FIFO_blk[8] = 1'b0;
    assign proc_3_TLF_FIFO_blk[8] = 1'b0;
    assign proc_3_input_sync_blk[8] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_3_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_3[8] = dl_detect_out ? proc_dep_vld_vec_3_reg[8] : (proc_3_data_FIFO_blk[8] | proc_3_data_PIPO_blk[8] | proc_3_start_FIFO_blk[8] | proc_3_TLF_FIFO_blk[8] | proc_3_input_sync_blk[8] | proc_3_output_sync_blk[8]);
    assign proc_3_data_FIFO_blk[9] = 1'b0;
    assign proc_3_data_PIPO_blk[9] = 1'b0;
    assign proc_3_start_FIFO_blk[9] = 1'b0;
    assign proc_3_TLF_FIFO_blk[9] = 1'b0;
    assign proc_3_input_sync_blk[9] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_3_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_3[9] = dl_detect_out ? proc_dep_vld_vec_3_reg[9] : (proc_3_data_FIFO_blk[9] | proc_3_data_PIPO_blk[9] | proc_3_start_FIFO_blk[9] | proc_3_TLF_FIFO_blk[9] | proc_3_input_sync_blk[9] | proc_3_output_sync_blk[9]);
    assign proc_3_data_FIFO_blk[10] = 1'b0;
    assign proc_3_data_PIPO_blk[10] = 1'b0;
    assign proc_3_start_FIFO_blk[10] = 1'b0;
    assign proc_3_TLF_FIFO_blk[10] = 1'b0;
    assign proc_3_input_sync_blk[10] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_3_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_3[10] = dl_detect_out ? proc_dep_vld_vec_3_reg[10] : (proc_3_data_FIFO_blk[10] | proc_3_data_PIPO_blk[10] | proc_3_start_FIFO_blk[10] | proc_3_TLF_FIFO_blk[10] | proc_3_input_sync_blk[10] | proc_3_output_sync_blk[10]);
    assign proc_3_data_FIFO_blk[11] = 1'b0;
    assign proc_3_data_PIPO_blk[11] = 1'b0;
    assign proc_3_start_FIFO_blk[11] = 1'b0;
    assign proc_3_TLF_FIFO_blk[11] = 1'b0;
    assign proc_3_input_sync_blk[11] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_3_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_3[11] = dl_detect_out ? proc_dep_vld_vec_3_reg[11] : (proc_3_data_FIFO_blk[11] | proc_3_data_PIPO_blk[11] | proc_3_start_FIFO_blk[11] | proc_3_TLF_FIFO_blk[11] | proc_3_input_sync_blk[11] | proc_3_output_sync_blk[11]);
    assign proc_3_data_FIFO_blk[12] = 1'b0;
    assign proc_3_data_PIPO_blk[12] = 1'b0;
    assign proc_3_start_FIFO_blk[12] = 1'b0;
    assign proc_3_TLF_FIFO_blk[12] = 1'b0;
    assign proc_3_input_sync_blk[12] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_3_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_3[12] = dl_detect_out ? proc_dep_vld_vec_3_reg[12] : (proc_3_data_FIFO_blk[12] | proc_3_data_PIPO_blk[12] | proc_3_start_FIFO_blk[12] | proc_3_TLF_FIFO_blk[12] | proc_3_input_sync_blk[12] | proc_3_output_sync_blk[12]);
    assign proc_3_data_FIFO_blk[13] = 1'b0;
    assign proc_3_data_PIPO_blk[13] = 1'b0;
    assign proc_3_start_FIFO_blk[13] = 1'b0;
    assign proc_3_TLF_FIFO_blk[13] = 1'b0;
    assign proc_3_input_sync_blk[13] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_3_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_3[13] = dl_detect_out ? proc_dep_vld_vec_3_reg[13] : (proc_3_data_FIFO_blk[13] | proc_3_data_PIPO_blk[13] | proc_3_start_FIFO_blk[13] | proc_3_TLF_FIFO_blk[13] | proc_3_input_sync_blk[13] | proc_3_output_sync_blk[13]);
    assign proc_3_data_FIFO_blk[14] = 1'b0;
    assign proc_3_data_PIPO_blk[14] = 1'b0;
    assign proc_3_start_FIFO_blk[14] = 1'b0;
    assign proc_3_TLF_FIFO_blk[14] = 1'b0;
    assign proc_3_input_sync_blk[14] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_3_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_3[14] = dl_detect_out ? proc_dep_vld_vec_3_reg[14] : (proc_3_data_FIFO_blk[14] | proc_3_data_PIPO_blk[14] | proc_3_start_FIFO_blk[14] | proc_3_TLF_FIFO_blk[14] | proc_3_input_sync_blk[14] | proc_3_output_sync_blk[14]);
    assign proc_3_data_FIFO_blk[15] = 1'b0;
    assign proc_3_data_PIPO_blk[15] = 1'b0;
    assign proc_3_start_FIFO_blk[15] = 1'b0;
    assign proc_3_TLF_FIFO_blk[15] = 1'b0;
    assign proc_3_input_sync_blk[15] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_3_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_3[15] = dl_detect_out ? proc_dep_vld_vec_3_reg[15] : (proc_3_data_FIFO_blk[15] | proc_3_data_PIPO_blk[15] | proc_3_start_FIFO_blk[15] | proc_3_TLF_FIFO_blk[15] | proc_3_input_sync_blk[15] | proc_3_output_sync_blk[15]);
    assign proc_3_data_FIFO_blk[16] = 1'b0;
    assign proc_3_data_PIPO_blk[16] = 1'b0;
    assign proc_3_start_FIFO_blk[16] = 1'b0;
    assign proc_3_TLF_FIFO_blk[16] = 1'b0;
    assign proc_3_input_sync_blk[16] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_3_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_3[16] = dl_detect_out ? proc_dep_vld_vec_3_reg[16] : (proc_3_data_FIFO_blk[16] | proc_3_data_PIPO_blk[16] | proc_3_start_FIFO_blk[16] | proc_3_TLF_FIFO_blk[16] | proc_3_input_sync_blk[16] | proc_3_output_sync_blk[16]);
    assign proc_3_data_FIFO_blk[17] = 1'b0;
    assign proc_3_data_PIPO_blk[17] = 1'b0;
    assign proc_3_start_FIFO_blk[17] = 1'b0;
    assign proc_3_TLF_FIFO_blk[17] = 1'b0;
    assign proc_3_input_sync_blk[17] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_3_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_3[17] = dl_detect_out ? proc_dep_vld_vec_3_reg[17] : (proc_3_data_FIFO_blk[17] | proc_3_data_PIPO_blk[17] | proc_3_start_FIFO_blk[17] | proc_3_TLF_FIFO_blk[17] | proc_3_input_sync_blk[17] | proc_3_output_sync_blk[17]);
    assign proc_3_data_FIFO_blk[18] = 1'b0;
    assign proc_3_data_PIPO_blk[18] = 1'b0;
    assign proc_3_start_FIFO_blk[18] = 1'b0;
    assign proc_3_TLF_FIFO_blk[18] = 1'b0;
    assign proc_3_input_sync_blk[18] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_3_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_3[18] = dl_detect_out ? proc_dep_vld_vec_3_reg[18] : (proc_3_data_FIFO_blk[18] | proc_3_data_PIPO_blk[18] | proc_3_start_FIFO_blk[18] | proc_3_TLF_FIFO_blk[18] | proc_3_input_sync_blk[18] | proc_3_output_sync_blk[18]);
    assign proc_3_data_FIFO_blk[19] = 1'b0;
    assign proc_3_data_PIPO_blk[19] = 1'b0;
    assign proc_3_start_FIFO_blk[19] = 1'b0;
    assign proc_3_TLF_FIFO_blk[19] = 1'b0;
    assign proc_3_input_sync_blk[19] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_3_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_3[19] = dl_detect_out ? proc_dep_vld_vec_3_reg[19] : (proc_3_data_FIFO_blk[19] | proc_3_data_PIPO_blk[19] | proc_3_start_FIFO_blk[19] | proc_3_TLF_FIFO_blk[19] | proc_3_input_sync_blk[19] | proc_3_output_sync_blk[19]);
    assign proc_3_data_FIFO_blk[20] = 1'b0;
    assign proc_3_data_PIPO_blk[20] = 1'b0;
    assign proc_3_start_FIFO_blk[20] = 1'b0;
    assign proc_3_TLF_FIFO_blk[20] = 1'b0;
    assign proc_3_input_sync_blk[20] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_3_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_3[20] = dl_detect_out ? proc_dep_vld_vec_3_reg[20] : (proc_3_data_FIFO_blk[20] | proc_3_data_PIPO_blk[20] | proc_3_start_FIFO_blk[20] | proc_3_TLF_FIFO_blk[20] | proc_3_input_sync_blk[20] | proc_3_output_sync_blk[20]);
    assign proc_3_data_FIFO_blk[21] = 1'b0;
    assign proc_3_data_PIPO_blk[21] = 1'b0;
    assign proc_3_start_FIFO_blk[21] = 1'b0;
    assign proc_3_TLF_FIFO_blk[21] = 1'b0;
    assign proc_3_input_sync_blk[21] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_3_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_3[21] = dl_detect_out ? proc_dep_vld_vec_3_reg[21] : (proc_3_data_FIFO_blk[21] | proc_3_data_PIPO_blk[21] | proc_3_start_FIFO_blk[21] | proc_3_TLF_FIFO_blk[21] | proc_3_input_sync_blk[21] | proc_3_output_sync_blk[21]);
    assign proc_3_data_FIFO_blk[22] = 1'b0;
    assign proc_3_data_PIPO_blk[22] = 1'b0;
    assign proc_3_start_FIFO_blk[22] = 1'b0;
    assign proc_3_TLF_FIFO_blk[22] = 1'b0;
    assign proc_3_input_sync_blk[22] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_3_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_3[22] = dl_detect_out ? proc_dep_vld_vec_3_reg[22] : (proc_3_data_FIFO_blk[22] | proc_3_data_PIPO_blk[22] | proc_3_start_FIFO_blk[22] | proc_3_TLF_FIFO_blk[22] | proc_3_input_sync_blk[22] | proc_3_output_sync_blk[22]);
    assign proc_3_data_FIFO_blk[23] = 1'b0;
    assign proc_3_data_PIPO_blk[23] = 1'b0;
    assign proc_3_start_FIFO_blk[23] = 1'b0;
    assign proc_3_TLF_FIFO_blk[23] = 1'b0;
    assign proc_3_input_sync_blk[23] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_3_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_3[23] = dl_detect_out ? proc_dep_vld_vec_3_reg[23] : (proc_3_data_FIFO_blk[23] | proc_3_data_PIPO_blk[23] | proc_3_start_FIFO_blk[23] | proc_3_TLF_FIFO_blk[23] | proc_3_input_sync_blk[23] | proc_3_output_sync_blk[23]);
    assign proc_3_data_FIFO_blk[24] = 1'b0;
    assign proc_3_data_PIPO_blk[24] = 1'b0;
    assign proc_3_start_FIFO_blk[24] = 1'b0;
    assign proc_3_TLF_FIFO_blk[24] = 1'b0;
    assign proc_3_input_sync_blk[24] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_3_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_3[24] = dl_detect_out ? proc_dep_vld_vec_3_reg[24] : (proc_3_data_FIFO_blk[24] | proc_3_data_PIPO_blk[24] | proc_3_start_FIFO_blk[24] | proc_3_TLF_FIFO_blk[24] | proc_3_input_sync_blk[24] | proc_3_output_sync_blk[24]);
    assign proc_3_data_FIFO_blk[25] = 1'b0;
    assign proc_3_data_PIPO_blk[25] = 1'b0;
    assign proc_3_start_FIFO_blk[25] = 1'b0;
    assign proc_3_TLF_FIFO_blk[25] = 1'b0;
    assign proc_3_input_sync_blk[25] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_3_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_3[25] = dl_detect_out ? proc_dep_vld_vec_3_reg[25] : (proc_3_data_FIFO_blk[25] | proc_3_data_PIPO_blk[25] | proc_3_start_FIFO_blk[25] | proc_3_TLF_FIFO_blk[25] | proc_3_input_sync_blk[25] | proc_3_output_sync_blk[25]);
    assign proc_3_data_FIFO_blk[26] = 1'b0;
    assign proc_3_data_PIPO_blk[26] = 1'b0;
    assign proc_3_start_FIFO_blk[26] = 1'b0;
    assign proc_3_TLF_FIFO_blk[26] = 1'b0;
    assign proc_3_input_sync_blk[26] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_3_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_3[26] = dl_detect_out ? proc_dep_vld_vec_3_reg[26] : (proc_3_data_FIFO_blk[26] | proc_3_data_PIPO_blk[26] | proc_3_start_FIFO_blk[26] | proc_3_TLF_FIFO_blk[26] | proc_3_input_sync_blk[26] | proc_3_output_sync_blk[26]);
    assign proc_3_data_FIFO_blk[27] = 1'b0;
    assign proc_3_data_PIPO_blk[27] = 1'b0;
    assign proc_3_start_FIFO_blk[27] = 1'b0;
    assign proc_3_TLF_FIFO_blk[27] = 1'b0;
    assign proc_3_input_sync_blk[27] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_3_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_3[27] = dl_detect_out ? proc_dep_vld_vec_3_reg[27] : (proc_3_data_FIFO_blk[27] | proc_3_data_PIPO_blk[27] | proc_3_start_FIFO_blk[27] | proc_3_TLF_FIFO_blk[27] | proc_3_input_sync_blk[27] | proc_3_output_sync_blk[27]);
    assign proc_3_data_FIFO_blk[28] = 1'b0;
    assign proc_3_data_PIPO_blk[28] = 1'b0;
    assign proc_3_start_FIFO_blk[28] = 1'b0;
    assign proc_3_TLF_FIFO_blk[28] = 1'b0;
    assign proc_3_input_sync_blk[28] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_3_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_3[28] = dl_detect_out ? proc_dep_vld_vec_3_reg[28] : (proc_3_data_FIFO_blk[28] | proc_3_data_PIPO_blk[28] | proc_3_start_FIFO_blk[28] | proc_3_TLF_FIFO_blk[28] | proc_3_input_sync_blk[28] | proc_3_output_sync_blk[28]);
    assign proc_3_data_FIFO_blk[29] = 1'b0;
    assign proc_3_data_PIPO_blk[29] = 1'b0;
    assign proc_3_start_FIFO_blk[29] = 1'b0;
    assign proc_3_TLF_FIFO_blk[29] = 1'b0;
    assign proc_3_input_sync_blk[29] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_3_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_3[29] = dl_detect_out ? proc_dep_vld_vec_3_reg[29] : (proc_3_data_FIFO_blk[29] | proc_3_data_PIPO_blk[29] | proc_3_start_FIFO_blk[29] | proc_3_TLF_FIFO_blk[29] | proc_3_input_sync_blk[29] | proc_3_output_sync_blk[29]);
    assign proc_3_data_FIFO_blk[30] = 1'b0;
    assign proc_3_data_PIPO_blk[30] = 1'b0;
    assign proc_3_start_FIFO_blk[30] = 1'b0;
    assign proc_3_TLF_FIFO_blk[30] = 1'b0;
    assign proc_3_input_sync_blk[30] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_3_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_3[30] = dl_detect_out ? proc_dep_vld_vec_3_reg[30] : (proc_3_data_FIFO_blk[30] | proc_3_data_PIPO_blk[30] | proc_3_start_FIFO_blk[30] | proc_3_TLF_FIFO_blk[30] | proc_3_input_sync_blk[30] | proc_3_output_sync_blk[30]);
    assign proc_3_data_FIFO_blk[31] = 1'b0;
    assign proc_3_data_PIPO_blk[31] = 1'b0;
    assign proc_3_start_FIFO_blk[31] = 1'b0;
    assign proc_3_TLF_FIFO_blk[31] = 1'b0;
    assign proc_3_input_sync_blk[31] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_3_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_3[31] = dl_detect_out ? proc_dep_vld_vec_3_reg[31] : (proc_3_data_FIFO_blk[31] | proc_3_data_PIPO_blk[31] | proc_3_start_FIFO_blk[31] | proc_3_TLF_FIFO_blk[31] | proc_3_input_sync_blk[31] | proc_3_output_sync_blk[31]);
    assign proc_3_data_FIFO_blk[32] = 1'b0;
    assign proc_3_data_PIPO_blk[32] = 1'b0;
    assign proc_3_start_FIFO_blk[32] = 1'b0;
    assign proc_3_TLF_FIFO_blk[32] = 1'b0;
    assign proc_3_input_sync_blk[32] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_3_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_3[32] = dl_detect_out ? proc_dep_vld_vec_3_reg[32] : (proc_3_data_FIFO_blk[32] | proc_3_data_PIPO_blk[32] | proc_3_start_FIFO_blk[32] | proc_3_TLF_FIFO_blk[32] | proc_3_input_sync_blk[32] | proc_3_output_sync_blk[32]);
    assign proc_3_data_FIFO_blk[33] = 1'b0;
    assign proc_3_data_PIPO_blk[33] = 1'b0;
    assign proc_3_start_FIFO_blk[33] = 1'b0;
    assign proc_3_TLF_FIFO_blk[33] = 1'b0;
    assign proc_3_input_sync_blk[33] = 1'b0 | (ap_sync_ReadB_U0_ap_ready & ReadB_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_3_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_3[33] = dl_detect_out ? proc_dep_vld_vec_3_reg[33] : (proc_3_data_FIFO_blk[33] | proc_3_data_PIPO_blk[33] | proc_3_start_FIFO_blk[33] | proc_3_TLF_FIFO_blk[33] | proc_3_input_sync_blk[33] | proc_3_output_sync_blk[33]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_3_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_3_reg <= proc_dep_vld_vec_3;
        end
    end
    assign in_chan_dep_vld_vec_3[0] = dep_chan_vld_0_3;
    assign in_chan_dep_data_vec_3[39 : 0] = dep_chan_data_0_3;
    assign token_in_vec_3[0] = token_0_3;
    assign in_chan_dep_vld_vec_3[1] = dep_chan_vld_1_3;
    assign in_chan_dep_data_vec_3[79 : 40] = dep_chan_data_1_3;
    assign token_in_vec_3[1] = token_1_3;
    assign in_chan_dep_vld_vec_3[2] = dep_chan_vld_4_3;
    assign in_chan_dep_data_vec_3[119 : 80] = dep_chan_data_4_3;
    assign token_in_vec_3[2] = token_4_3;
    assign in_chan_dep_vld_vec_3[3] = dep_chan_vld_6_3;
    assign in_chan_dep_data_vec_3[159 : 120] = dep_chan_data_6_3;
    assign token_in_vec_3[3] = token_6_3;
    assign in_chan_dep_vld_vec_3[4] = dep_chan_vld_7_3;
    assign in_chan_dep_data_vec_3[199 : 160] = dep_chan_data_7_3;
    assign token_in_vec_3[4] = token_7_3;
    assign in_chan_dep_vld_vec_3[5] = dep_chan_vld_8_3;
    assign in_chan_dep_data_vec_3[239 : 200] = dep_chan_data_8_3;
    assign token_in_vec_3[5] = token_8_3;
    assign in_chan_dep_vld_vec_3[6] = dep_chan_vld_9_3;
    assign in_chan_dep_data_vec_3[279 : 240] = dep_chan_data_9_3;
    assign token_in_vec_3[6] = token_9_3;
    assign in_chan_dep_vld_vec_3[7] = dep_chan_vld_10_3;
    assign in_chan_dep_data_vec_3[319 : 280] = dep_chan_data_10_3;
    assign token_in_vec_3[7] = token_10_3;
    assign in_chan_dep_vld_vec_3[8] = dep_chan_vld_11_3;
    assign in_chan_dep_data_vec_3[359 : 320] = dep_chan_data_11_3;
    assign token_in_vec_3[8] = token_11_3;
    assign in_chan_dep_vld_vec_3[9] = dep_chan_vld_12_3;
    assign in_chan_dep_data_vec_3[399 : 360] = dep_chan_data_12_3;
    assign token_in_vec_3[9] = token_12_3;
    assign in_chan_dep_vld_vec_3[10] = dep_chan_vld_13_3;
    assign in_chan_dep_data_vec_3[439 : 400] = dep_chan_data_13_3;
    assign token_in_vec_3[10] = token_13_3;
    assign in_chan_dep_vld_vec_3[11] = dep_chan_vld_14_3;
    assign in_chan_dep_data_vec_3[479 : 440] = dep_chan_data_14_3;
    assign token_in_vec_3[11] = token_14_3;
    assign in_chan_dep_vld_vec_3[12] = dep_chan_vld_15_3;
    assign in_chan_dep_data_vec_3[519 : 480] = dep_chan_data_15_3;
    assign token_in_vec_3[12] = token_15_3;
    assign in_chan_dep_vld_vec_3[13] = dep_chan_vld_16_3;
    assign in_chan_dep_data_vec_3[559 : 520] = dep_chan_data_16_3;
    assign token_in_vec_3[13] = token_16_3;
    assign in_chan_dep_vld_vec_3[14] = dep_chan_vld_17_3;
    assign in_chan_dep_data_vec_3[599 : 560] = dep_chan_data_17_3;
    assign token_in_vec_3[14] = token_17_3;
    assign in_chan_dep_vld_vec_3[15] = dep_chan_vld_18_3;
    assign in_chan_dep_data_vec_3[639 : 600] = dep_chan_data_18_3;
    assign token_in_vec_3[15] = token_18_3;
    assign in_chan_dep_vld_vec_3[16] = dep_chan_vld_19_3;
    assign in_chan_dep_data_vec_3[679 : 640] = dep_chan_data_19_3;
    assign token_in_vec_3[16] = token_19_3;
    assign in_chan_dep_vld_vec_3[17] = dep_chan_vld_20_3;
    assign in_chan_dep_data_vec_3[719 : 680] = dep_chan_data_20_3;
    assign token_in_vec_3[17] = token_20_3;
    assign in_chan_dep_vld_vec_3[18] = dep_chan_vld_21_3;
    assign in_chan_dep_data_vec_3[759 : 720] = dep_chan_data_21_3;
    assign token_in_vec_3[18] = token_21_3;
    assign in_chan_dep_vld_vec_3[19] = dep_chan_vld_22_3;
    assign in_chan_dep_data_vec_3[799 : 760] = dep_chan_data_22_3;
    assign token_in_vec_3[19] = token_22_3;
    assign in_chan_dep_vld_vec_3[20] = dep_chan_vld_23_3;
    assign in_chan_dep_data_vec_3[839 : 800] = dep_chan_data_23_3;
    assign token_in_vec_3[20] = token_23_3;
    assign in_chan_dep_vld_vec_3[21] = dep_chan_vld_24_3;
    assign in_chan_dep_data_vec_3[879 : 840] = dep_chan_data_24_3;
    assign token_in_vec_3[21] = token_24_3;
    assign in_chan_dep_vld_vec_3[22] = dep_chan_vld_25_3;
    assign in_chan_dep_data_vec_3[919 : 880] = dep_chan_data_25_3;
    assign token_in_vec_3[22] = token_25_3;
    assign in_chan_dep_vld_vec_3[23] = dep_chan_vld_26_3;
    assign in_chan_dep_data_vec_3[959 : 920] = dep_chan_data_26_3;
    assign token_in_vec_3[23] = token_26_3;
    assign in_chan_dep_vld_vec_3[24] = dep_chan_vld_27_3;
    assign in_chan_dep_data_vec_3[999 : 960] = dep_chan_data_27_3;
    assign token_in_vec_3[24] = token_27_3;
    assign in_chan_dep_vld_vec_3[25] = dep_chan_vld_28_3;
    assign in_chan_dep_data_vec_3[1039 : 1000] = dep_chan_data_28_3;
    assign token_in_vec_3[25] = token_28_3;
    assign in_chan_dep_vld_vec_3[26] = dep_chan_vld_29_3;
    assign in_chan_dep_data_vec_3[1079 : 1040] = dep_chan_data_29_3;
    assign token_in_vec_3[26] = token_29_3;
    assign in_chan_dep_vld_vec_3[27] = dep_chan_vld_30_3;
    assign in_chan_dep_data_vec_3[1119 : 1080] = dep_chan_data_30_3;
    assign token_in_vec_3[27] = token_30_3;
    assign in_chan_dep_vld_vec_3[28] = dep_chan_vld_31_3;
    assign in_chan_dep_data_vec_3[1159 : 1120] = dep_chan_data_31_3;
    assign token_in_vec_3[28] = token_31_3;
    assign in_chan_dep_vld_vec_3[29] = dep_chan_vld_32_3;
    assign in_chan_dep_data_vec_3[1199 : 1160] = dep_chan_data_32_3;
    assign token_in_vec_3[29] = token_32_3;
    assign in_chan_dep_vld_vec_3[30] = dep_chan_vld_33_3;
    assign in_chan_dep_data_vec_3[1239 : 1200] = dep_chan_data_33_3;
    assign token_in_vec_3[30] = token_33_3;
    assign in_chan_dep_vld_vec_3[31] = dep_chan_vld_34_3;
    assign in_chan_dep_data_vec_3[1279 : 1240] = dep_chan_data_34_3;
    assign token_in_vec_3[31] = token_34_3;
    assign in_chan_dep_vld_vec_3[32] = dep_chan_vld_35_3;
    assign in_chan_dep_data_vec_3[1319 : 1280] = dep_chan_data_35_3;
    assign token_in_vec_3[32] = token_35_3;
    assign in_chan_dep_vld_vec_3[33] = dep_chan_vld_36_3;
    assign in_chan_dep_data_vec_3[1359 : 1320] = dep_chan_data_36_3;
    assign token_in_vec_3[33] = token_36_3;
    assign dep_chan_vld_3_4 = out_chan_dep_vld_vec_3[0];
    assign dep_chan_data_3_4 = out_chan_dep_data_3;
    assign token_3_4 = token_out_vec_3[0];
    assign dep_chan_vld_3_0 = out_chan_dep_vld_vec_3[1];
    assign dep_chan_data_3_0 = out_chan_dep_data_3;
    assign token_3_0 = token_out_vec_3[1];
    assign dep_chan_vld_3_1 = out_chan_dep_vld_vec_3[2];
    assign dep_chan_data_3_1 = out_chan_dep_data_3;
    assign token_3_1 = token_out_vec_3[2];
    assign dep_chan_vld_3_6 = out_chan_dep_vld_vec_3[3];
    assign dep_chan_data_3_6 = out_chan_dep_data_3;
    assign token_3_6 = token_out_vec_3[3];
    assign dep_chan_vld_3_7 = out_chan_dep_vld_vec_3[4];
    assign dep_chan_data_3_7 = out_chan_dep_data_3;
    assign token_3_7 = token_out_vec_3[4];
    assign dep_chan_vld_3_8 = out_chan_dep_vld_vec_3[5];
    assign dep_chan_data_3_8 = out_chan_dep_data_3;
    assign token_3_8 = token_out_vec_3[5];
    assign dep_chan_vld_3_9 = out_chan_dep_vld_vec_3[6];
    assign dep_chan_data_3_9 = out_chan_dep_data_3;
    assign token_3_9 = token_out_vec_3[6];
    assign dep_chan_vld_3_10 = out_chan_dep_vld_vec_3[7];
    assign dep_chan_data_3_10 = out_chan_dep_data_3;
    assign token_3_10 = token_out_vec_3[7];
    assign dep_chan_vld_3_11 = out_chan_dep_vld_vec_3[8];
    assign dep_chan_data_3_11 = out_chan_dep_data_3;
    assign token_3_11 = token_out_vec_3[8];
    assign dep_chan_vld_3_12 = out_chan_dep_vld_vec_3[9];
    assign dep_chan_data_3_12 = out_chan_dep_data_3;
    assign token_3_12 = token_out_vec_3[9];
    assign dep_chan_vld_3_13 = out_chan_dep_vld_vec_3[10];
    assign dep_chan_data_3_13 = out_chan_dep_data_3;
    assign token_3_13 = token_out_vec_3[10];
    assign dep_chan_vld_3_14 = out_chan_dep_vld_vec_3[11];
    assign dep_chan_data_3_14 = out_chan_dep_data_3;
    assign token_3_14 = token_out_vec_3[11];
    assign dep_chan_vld_3_15 = out_chan_dep_vld_vec_3[12];
    assign dep_chan_data_3_15 = out_chan_dep_data_3;
    assign token_3_15 = token_out_vec_3[12];
    assign dep_chan_vld_3_16 = out_chan_dep_vld_vec_3[13];
    assign dep_chan_data_3_16 = out_chan_dep_data_3;
    assign token_3_16 = token_out_vec_3[13];
    assign dep_chan_vld_3_17 = out_chan_dep_vld_vec_3[14];
    assign dep_chan_data_3_17 = out_chan_dep_data_3;
    assign token_3_17 = token_out_vec_3[14];
    assign dep_chan_vld_3_18 = out_chan_dep_vld_vec_3[15];
    assign dep_chan_data_3_18 = out_chan_dep_data_3;
    assign token_3_18 = token_out_vec_3[15];
    assign dep_chan_vld_3_19 = out_chan_dep_vld_vec_3[16];
    assign dep_chan_data_3_19 = out_chan_dep_data_3;
    assign token_3_19 = token_out_vec_3[16];
    assign dep_chan_vld_3_20 = out_chan_dep_vld_vec_3[17];
    assign dep_chan_data_3_20 = out_chan_dep_data_3;
    assign token_3_20 = token_out_vec_3[17];
    assign dep_chan_vld_3_21 = out_chan_dep_vld_vec_3[18];
    assign dep_chan_data_3_21 = out_chan_dep_data_3;
    assign token_3_21 = token_out_vec_3[18];
    assign dep_chan_vld_3_22 = out_chan_dep_vld_vec_3[19];
    assign dep_chan_data_3_22 = out_chan_dep_data_3;
    assign token_3_22 = token_out_vec_3[19];
    assign dep_chan_vld_3_23 = out_chan_dep_vld_vec_3[20];
    assign dep_chan_data_3_23 = out_chan_dep_data_3;
    assign token_3_23 = token_out_vec_3[20];
    assign dep_chan_vld_3_24 = out_chan_dep_vld_vec_3[21];
    assign dep_chan_data_3_24 = out_chan_dep_data_3;
    assign token_3_24 = token_out_vec_3[21];
    assign dep_chan_vld_3_25 = out_chan_dep_vld_vec_3[22];
    assign dep_chan_data_3_25 = out_chan_dep_data_3;
    assign token_3_25 = token_out_vec_3[22];
    assign dep_chan_vld_3_26 = out_chan_dep_vld_vec_3[23];
    assign dep_chan_data_3_26 = out_chan_dep_data_3;
    assign token_3_26 = token_out_vec_3[23];
    assign dep_chan_vld_3_27 = out_chan_dep_vld_vec_3[24];
    assign dep_chan_data_3_27 = out_chan_dep_data_3;
    assign token_3_27 = token_out_vec_3[24];
    assign dep_chan_vld_3_28 = out_chan_dep_vld_vec_3[25];
    assign dep_chan_data_3_28 = out_chan_dep_data_3;
    assign token_3_28 = token_out_vec_3[25];
    assign dep_chan_vld_3_29 = out_chan_dep_vld_vec_3[26];
    assign dep_chan_data_3_29 = out_chan_dep_data_3;
    assign token_3_29 = token_out_vec_3[26];
    assign dep_chan_vld_3_30 = out_chan_dep_vld_vec_3[27];
    assign dep_chan_data_3_30 = out_chan_dep_data_3;
    assign token_3_30 = token_out_vec_3[27];
    assign dep_chan_vld_3_31 = out_chan_dep_vld_vec_3[28];
    assign dep_chan_data_3_31 = out_chan_dep_data_3;
    assign token_3_31 = token_out_vec_3[28];
    assign dep_chan_vld_3_32 = out_chan_dep_vld_vec_3[29];
    assign dep_chan_data_3_32 = out_chan_dep_data_3;
    assign token_3_32 = token_out_vec_3[29];
    assign dep_chan_vld_3_33 = out_chan_dep_vld_vec_3[30];
    assign dep_chan_data_3_33 = out_chan_dep_data_3;
    assign token_3_33 = token_out_vec_3[30];
    assign dep_chan_vld_3_34 = out_chan_dep_vld_vec_3[31];
    assign dep_chan_data_3_34 = out_chan_dep_data_3;
    assign token_3_34 = token_out_vec_3[31];
    assign dep_chan_vld_3_35 = out_chan_dep_vld_vec_3[32];
    assign dep_chan_data_3_35 = out_chan_dep_data_3;
    assign token_3_35 = token_out_vec_3[32];
    assign dep_chan_vld_3_36 = out_chan_dep_vld_vec_3[33];
    assign dep_chan_data_3_36 = out_chan_dep_data_3;
    assign token_3_36 = token_out_vec_3[33];

    // Process: ConvertWidthB_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 4, 2, 2) MatrixMultiplicationKernel_hls_deadlock_detect_unit_4 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_4),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_4),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_4),
        .token_in_vec(token_in_vec_4),
        .dl_detect_in(dl_detect_out),
        .origin(origin[4]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_4),
        .out_chan_dep_data(out_chan_dep_data_4),
        .token_out_vec(token_out_vec_4),
        .dl_detect_out(dl_in_vec[4]));

    assign proc_4_data_FIFO_blk[0] = 1'b0 | (~ConvertWidthB_U0.grp_ConvertWidthB_Pipeline_ConvertWidthB_Outer_ConvertWidthB_Memory_fu_98.bMemory_blk_n) | (~ConvertWidthB_U0.size_n_blk_n) | (~ConvertWidthB_U0.size_k_blk_n) | (~ConvertWidthB_U0.size_m_blk_n);
    assign proc_4_data_PIPO_blk[0] = 1'b0;
    assign proc_4_start_FIFO_blk[0] = 1'b0 | (~start_for_ConvertWidthB_U0_U.if_empty_n & ConvertWidthB_U0.ap_idle & ~start_for_ConvertWidthB_U0_U.if_write);
    assign proc_4_TLF_FIFO_blk[0] = 1'b0;
    assign proc_4_input_sync_blk[0] = 1'b0;
    assign proc_4_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_4[0] = dl_detect_out ? proc_dep_vld_vec_4_reg[0] : (proc_4_data_FIFO_blk[0] | proc_4_data_PIPO_blk[0] | proc_4_start_FIFO_blk[0] | proc_4_TLF_FIFO_blk[0] | proc_4_input_sync_blk[0] | proc_4_output_sync_blk[0]);
    assign proc_4_data_FIFO_blk[1] = 1'b0 | (~ConvertWidthB_U0.grp_ConvertWidthB_Pipeline_ConvertWidthB_Outer_ConvertWidthB_Memory_fu_98.bFeed_blk_n) | (~ConvertWidthB_U0.size_n_c3_blk_n) | (~ConvertWidthB_U0.size_k_c6_blk_n) | (~ConvertWidthB_U0.size_m_c11_blk_n);
    assign proc_4_data_PIPO_blk[1] = 1'b0;
    assign proc_4_start_FIFO_blk[1] = 1'b0 | (~start_for_FeedB_U0_U.if_full_n & ConvertWidthB_U0.ap_start & ~ConvertWidthB_U0.real_start & (trans_in_cnt_2 == trans_out_cnt_2) & ~start_for_FeedB_U0_U.if_read);
    assign proc_4_TLF_FIFO_blk[1] = 1'b0;
    assign proc_4_input_sync_blk[1] = 1'b0;
    assign proc_4_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_4[1] = dl_detect_out ? proc_dep_vld_vec_4_reg[1] : (proc_4_data_FIFO_blk[1] | proc_4_data_PIPO_blk[1] | proc_4_start_FIFO_blk[1] | proc_4_TLF_FIFO_blk[1] | proc_4_input_sync_blk[1] | proc_4_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_4_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_4_reg <= proc_dep_vld_vec_4;
        end
    end
    assign in_chan_dep_vld_vec_4[0] = dep_chan_vld_3_4;
    assign in_chan_dep_data_vec_4[39 : 0] = dep_chan_data_3_4;
    assign token_in_vec_4[0] = token_3_4;
    assign in_chan_dep_vld_vec_4[1] = dep_chan_vld_5_4;
    assign in_chan_dep_data_vec_4[79 : 40] = dep_chan_data_5_4;
    assign token_in_vec_4[1] = token_5_4;
    assign dep_chan_vld_4_3 = out_chan_dep_vld_vec_4[0];
    assign dep_chan_data_4_3 = out_chan_dep_data_4;
    assign token_4_3 = token_out_vec_4[0];
    assign dep_chan_vld_4_5 = out_chan_dep_vld_vec_4[1];
    assign dep_chan_data_4_5 = out_chan_dep_data_4;
    assign token_4_5 = token_out_vec_4[1];

    // Process: FeedB_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 5, 2, 2) MatrixMultiplicationKernel_hls_deadlock_detect_unit_5 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_5),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_5),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_5),
        .token_in_vec(token_in_vec_5),
        .dl_detect_in(dl_detect_out),
        .origin(origin[5]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_5),
        .out_chan_dep_data(out_chan_dep_data_5),
        .token_out_vec(token_out_vec_5),
        .dl_detect_out(dl_in_vec[5]));

    assign proc_5_data_FIFO_blk[0] = 1'b0 | (~FeedB_U0.grp_FeedB_Pipeline_FeedB_Pipeline_N_FeedB_Pipeline_M_fu_123.bFeed_blk_n) | (~FeedB_U0.size_n_blk_n) | (~FeedB_U0.size_k_blk_n) | (~FeedB_U0.size_m_blk_n);
    assign proc_5_data_PIPO_blk[0] = 1'b0;
    assign proc_5_start_FIFO_blk[0] = 1'b0 | (~start_for_FeedB_U0_U.if_empty_n & FeedB_U0.ap_idle & ~start_for_FeedB_U0_U.if_write);
    assign proc_5_TLF_FIFO_blk[0] = 1'b0;
    assign proc_5_input_sync_blk[0] = 1'b0;
    assign proc_5_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_5[0] = dl_detect_out ? proc_dep_vld_vec_5_reg[0] : (proc_5_data_FIFO_blk[0] | proc_5_data_PIPO_blk[0] | proc_5_start_FIFO_blk[0] | proc_5_TLF_FIFO_blk[0] | proc_5_input_sync_blk[0] | proc_5_output_sync_blk[0]);
    assign proc_5_data_FIFO_blk[1] = 1'b0 | (~FeedB_U0.grp_FeedB_Pipeline_FeedB_Pipeline_N_FeedB_Pipeline_M_fu_123.bPipes_0_blk_n);
    assign proc_5_data_PIPO_blk[1] = 1'b0;
    assign proc_5_start_FIFO_blk[1] = 1'b0;
    assign proc_5_TLF_FIFO_blk[1] = 1'b0;
    assign proc_5_input_sync_blk[1] = 1'b0;
    assign proc_5_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_5[1] = dl_detect_out ? proc_dep_vld_vec_5_reg[1] : (proc_5_data_FIFO_blk[1] | proc_5_data_PIPO_blk[1] | proc_5_start_FIFO_blk[1] | proc_5_TLF_FIFO_blk[1] | proc_5_input_sync_blk[1] | proc_5_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_5_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_5_reg <= proc_dep_vld_vec_5;
        end
    end
    assign in_chan_dep_vld_vec_5[0] = dep_chan_vld_4_5;
    assign in_chan_dep_data_vec_5[39 : 0] = dep_chan_data_4_5;
    assign token_in_vec_5[0] = token_4_5;
    assign in_chan_dep_vld_vec_5[1] = dep_chan_vld_6_5;
    assign in_chan_dep_data_vec_5[79 : 40] = dep_chan_data_6_5;
    assign token_in_vec_5[1] = token_6_5;
    assign dep_chan_vld_5_4 = out_chan_dep_vld_vec_5[0];
    assign dep_chan_data_5_4 = out_chan_dep_data_5;
    assign token_5_4 = token_out_vec_5[0];
    assign dep_chan_vld_5_6 = out_chan_dep_vld_vec_5[1];
    assign dep_chan_data_5_6 = out_chan_dep_data_5;
    assign token_5_6 = token_out_vec_5[1];

    // Process: ProcessingElement_1_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 6, 36, 36) MatrixMultiplicationKernel_hls_deadlock_detect_unit_6 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_6),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_6),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_6),
        .token_in_vec(token_in_vec_6),
        .dl_detect_in(dl_detect_out),
        .origin(origin[6]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_6),
        .out_chan_dep_data(out_chan_dep_data_6),
        .token_out_vec(token_out_vec_6),
        .dl_detect_out(dl_in_vec[6]));

    assign proc_6_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_Pipeline_N_Pipeline_M_fu_189.aPipes_0_blk_n);
    assign proc_6_data_PIPO_blk[0] = 1'b0;
    assign proc_6_start_FIFO_blk[0] = 1'b0;
    assign proc_6_TLF_FIFO_blk[0] = 1'b0;
    assign proc_6_input_sync_blk[0] = 1'b0;
    assign proc_6_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_6[0] = dl_detect_out ? proc_dep_vld_vec_6_reg[0] : (proc_6_data_FIFO_blk[0] | proc_6_data_PIPO_blk[0] | proc_6_start_FIFO_blk[0] | proc_6_TLF_FIFO_blk[0] | proc_6_input_sync_blk[0] | proc_6_output_sync_blk[0]);
    assign proc_6_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_Pipeline_N_Pipeline_M_fu_189.aPipes_1_blk_n) | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_Pipeline_N_Pipeline_M_fu_189.bPipes_1_blk_n) | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_WriteC_Flattened_fu_211.cPipes_1_blk_n);
    assign proc_6_data_PIPO_blk[1] = 1'b0;
    assign proc_6_start_FIFO_blk[1] = 1'b0;
    assign proc_6_TLF_FIFO_blk[1] = 1'b0;
    assign proc_6_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_6_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_6[1] = dl_detect_out ? proc_dep_vld_vec_6_reg[1] : (proc_6_data_FIFO_blk[1] | proc_6_data_PIPO_blk[1] | proc_6_start_FIFO_blk[1] | proc_6_TLF_FIFO_blk[1] | proc_6_input_sync_blk[1] | proc_6_output_sync_blk[1]);
    assign proc_6_data_FIFO_blk[2] = 1'b0 | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_Pipeline_N_Pipeline_M_fu_189.bPipes_0_blk_n);
    assign proc_6_data_PIPO_blk[2] = 1'b0;
    assign proc_6_start_FIFO_blk[2] = 1'b0;
    assign proc_6_TLF_FIFO_blk[2] = 1'b0;
    assign proc_6_input_sync_blk[2] = 1'b0;
    assign proc_6_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_6[2] = dl_detect_out ? proc_dep_vld_vec_6_reg[2] : (proc_6_data_FIFO_blk[2] | proc_6_data_PIPO_blk[2] | proc_6_start_FIFO_blk[2] | proc_6_TLF_FIFO_blk[2] | proc_6_input_sync_blk[2] | proc_6_output_sync_blk[2]);
    assign proc_6_data_FIFO_blk[3] = 1'b0 | (~ProcessingElement_1_U0.grp_ProcessingElement_1_Pipeline_WriteC_Flattened_fu_211.cPipes_0_blk_n) | (~ProcessingElement_1_U0.size_n_c1_blk_n) | (~ProcessingElement_1_U0.size_m_c9_blk_n);
    assign proc_6_data_PIPO_blk[3] = 1'b0;
    assign proc_6_start_FIFO_blk[3] = 1'b0 | (~start_for_ConvertWidthC_U0_U.if_full_n & ProcessingElement_1_U0.ap_start & ~ProcessingElement_1_U0.real_start & (trans_in_cnt_4 == trans_out_cnt_4) & ~start_for_ConvertWidthC_U0_U.if_read);
    assign proc_6_TLF_FIFO_blk[3] = 1'b0;
    assign proc_6_input_sync_blk[3] = 1'b0;
    assign proc_6_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_6[3] = dl_detect_out ? proc_dep_vld_vec_6_reg[3] : (proc_6_data_FIFO_blk[3] | proc_6_data_PIPO_blk[3] | proc_6_start_FIFO_blk[3] | proc_6_TLF_FIFO_blk[3] | proc_6_input_sync_blk[3] | proc_6_output_sync_blk[3]);
    assign proc_6_data_FIFO_blk[4] = 1'b0;
    assign proc_6_data_PIPO_blk[4] = 1'b0;
    assign proc_6_start_FIFO_blk[4] = 1'b0;
    assign proc_6_TLF_FIFO_blk[4] = 1'b0;
    assign proc_6_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_6_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_6[4] = dl_detect_out ? proc_dep_vld_vec_6_reg[4] : (proc_6_data_FIFO_blk[4] | proc_6_data_PIPO_blk[4] | proc_6_start_FIFO_blk[4] | proc_6_TLF_FIFO_blk[4] | proc_6_input_sync_blk[4] | proc_6_output_sync_blk[4]);
    assign proc_6_data_FIFO_blk[5] = 1'b0;
    assign proc_6_data_PIPO_blk[5] = 1'b0;
    assign proc_6_start_FIFO_blk[5] = 1'b0;
    assign proc_6_TLF_FIFO_blk[5] = 1'b0;
    assign proc_6_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_6_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_6[5] = dl_detect_out ? proc_dep_vld_vec_6_reg[5] : (proc_6_data_FIFO_blk[5] | proc_6_data_PIPO_blk[5] | proc_6_start_FIFO_blk[5] | proc_6_TLF_FIFO_blk[5] | proc_6_input_sync_blk[5] | proc_6_output_sync_blk[5]);
    assign proc_6_data_FIFO_blk[6] = 1'b0;
    assign proc_6_data_PIPO_blk[6] = 1'b0;
    assign proc_6_start_FIFO_blk[6] = 1'b0;
    assign proc_6_TLF_FIFO_blk[6] = 1'b0;
    assign proc_6_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_6_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_6[6] = dl_detect_out ? proc_dep_vld_vec_6_reg[6] : (proc_6_data_FIFO_blk[6] | proc_6_data_PIPO_blk[6] | proc_6_start_FIFO_blk[6] | proc_6_TLF_FIFO_blk[6] | proc_6_input_sync_blk[6] | proc_6_output_sync_blk[6]);
    assign proc_6_data_FIFO_blk[7] = 1'b0;
    assign proc_6_data_PIPO_blk[7] = 1'b0;
    assign proc_6_start_FIFO_blk[7] = 1'b0;
    assign proc_6_TLF_FIFO_blk[7] = 1'b0;
    assign proc_6_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_6_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_6[7] = dl_detect_out ? proc_dep_vld_vec_6_reg[7] : (proc_6_data_FIFO_blk[7] | proc_6_data_PIPO_blk[7] | proc_6_start_FIFO_blk[7] | proc_6_TLF_FIFO_blk[7] | proc_6_input_sync_blk[7] | proc_6_output_sync_blk[7]);
    assign proc_6_data_FIFO_blk[8] = 1'b0;
    assign proc_6_data_PIPO_blk[8] = 1'b0;
    assign proc_6_start_FIFO_blk[8] = 1'b0;
    assign proc_6_TLF_FIFO_blk[8] = 1'b0;
    assign proc_6_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_6_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_6[8] = dl_detect_out ? proc_dep_vld_vec_6_reg[8] : (proc_6_data_FIFO_blk[8] | proc_6_data_PIPO_blk[8] | proc_6_start_FIFO_blk[8] | proc_6_TLF_FIFO_blk[8] | proc_6_input_sync_blk[8] | proc_6_output_sync_blk[8]);
    assign proc_6_data_FIFO_blk[9] = 1'b0;
    assign proc_6_data_PIPO_blk[9] = 1'b0;
    assign proc_6_start_FIFO_blk[9] = 1'b0;
    assign proc_6_TLF_FIFO_blk[9] = 1'b0;
    assign proc_6_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_6_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_6[9] = dl_detect_out ? proc_dep_vld_vec_6_reg[9] : (proc_6_data_FIFO_blk[9] | proc_6_data_PIPO_blk[9] | proc_6_start_FIFO_blk[9] | proc_6_TLF_FIFO_blk[9] | proc_6_input_sync_blk[9] | proc_6_output_sync_blk[9]);
    assign proc_6_data_FIFO_blk[10] = 1'b0;
    assign proc_6_data_PIPO_blk[10] = 1'b0;
    assign proc_6_start_FIFO_blk[10] = 1'b0;
    assign proc_6_TLF_FIFO_blk[10] = 1'b0;
    assign proc_6_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_6_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_6[10] = dl_detect_out ? proc_dep_vld_vec_6_reg[10] : (proc_6_data_FIFO_blk[10] | proc_6_data_PIPO_blk[10] | proc_6_start_FIFO_blk[10] | proc_6_TLF_FIFO_blk[10] | proc_6_input_sync_blk[10] | proc_6_output_sync_blk[10]);
    assign proc_6_data_FIFO_blk[11] = 1'b0;
    assign proc_6_data_PIPO_blk[11] = 1'b0;
    assign proc_6_start_FIFO_blk[11] = 1'b0;
    assign proc_6_TLF_FIFO_blk[11] = 1'b0;
    assign proc_6_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_6_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_6[11] = dl_detect_out ? proc_dep_vld_vec_6_reg[11] : (proc_6_data_FIFO_blk[11] | proc_6_data_PIPO_blk[11] | proc_6_start_FIFO_blk[11] | proc_6_TLF_FIFO_blk[11] | proc_6_input_sync_blk[11] | proc_6_output_sync_blk[11]);
    assign proc_6_data_FIFO_blk[12] = 1'b0;
    assign proc_6_data_PIPO_blk[12] = 1'b0;
    assign proc_6_start_FIFO_blk[12] = 1'b0;
    assign proc_6_TLF_FIFO_blk[12] = 1'b0;
    assign proc_6_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_6_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_6[12] = dl_detect_out ? proc_dep_vld_vec_6_reg[12] : (proc_6_data_FIFO_blk[12] | proc_6_data_PIPO_blk[12] | proc_6_start_FIFO_blk[12] | proc_6_TLF_FIFO_blk[12] | proc_6_input_sync_blk[12] | proc_6_output_sync_blk[12]);
    assign proc_6_data_FIFO_blk[13] = 1'b0;
    assign proc_6_data_PIPO_blk[13] = 1'b0;
    assign proc_6_start_FIFO_blk[13] = 1'b0;
    assign proc_6_TLF_FIFO_blk[13] = 1'b0;
    assign proc_6_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_6_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_6[13] = dl_detect_out ? proc_dep_vld_vec_6_reg[13] : (proc_6_data_FIFO_blk[13] | proc_6_data_PIPO_blk[13] | proc_6_start_FIFO_blk[13] | proc_6_TLF_FIFO_blk[13] | proc_6_input_sync_blk[13] | proc_6_output_sync_blk[13]);
    assign proc_6_data_FIFO_blk[14] = 1'b0;
    assign proc_6_data_PIPO_blk[14] = 1'b0;
    assign proc_6_start_FIFO_blk[14] = 1'b0;
    assign proc_6_TLF_FIFO_blk[14] = 1'b0;
    assign proc_6_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_6_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_6[14] = dl_detect_out ? proc_dep_vld_vec_6_reg[14] : (proc_6_data_FIFO_blk[14] | proc_6_data_PIPO_blk[14] | proc_6_start_FIFO_blk[14] | proc_6_TLF_FIFO_blk[14] | proc_6_input_sync_blk[14] | proc_6_output_sync_blk[14]);
    assign proc_6_data_FIFO_blk[15] = 1'b0;
    assign proc_6_data_PIPO_blk[15] = 1'b0;
    assign proc_6_start_FIFO_blk[15] = 1'b0;
    assign proc_6_TLF_FIFO_blk[15] = 1'b0;
    assign proc_6_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_6_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_6[15] = dl_detect_out ? proc_dep_vld_vec_6_reg[15] : (proc_6_data_FIFO_blk[15] | proc_6_data_PIPO_blk[15] | proc_6_start_FIFO_blk[15] | proc_6_TLF_FIFO_blk[15] | proc_6_input_sync_blk[15] | proc_6_output_sync_blk[15]);
    assign proc_6_data_FIFO_blk[16] = 1'b0;
    assign proc_6_data_PIPO_blk[16] = 1'b0;
    assign proc_6_start_FIFO_blk[16] = 1'b0;
    assign proc_6_TLF_FIFO_blk[16] = 1'b0;
    assign proc_6_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_6_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_6[16] = dl_detect_out ? proc_dep_vld_vec_6_reg[16] : (proc_6_data_FIFO_blk[16] | proc_6_data_PIPO_blk[16] | proc_6_start_FIFO_blk[16] | proc_6_TLF_FIFO_blk[16] | proc_6_input_sync_blk[16] | proc_6_output_sync_blk[16]);
    assign proc_6_data_FIFO_blk[17] = 1'b0;
    assign proc_6_data_PIPO_blk[17] = 1'b0;
    assign proc_6_start_FIFO_blk[17] = 1'b0;
    assign proc_6_TLF_FIFO_blk[17] = 1'b0;
    assign proc_6_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_6_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_6[17] = dl_detect_out ? proc_dep_vld_vec_6_reg[17] : (proc_6_data_FIFO_blk[17] | proc_6_data_PIPO_blk[17] | proc_6_start_FIFO_blk[17] | proc_6_TLF_FIFO_blk[17] | proc_6_input_sync_blk[17] | proc_6_output_sync_blk[17]);
    assign proc_6_data_FIFO_blk[18] = 1'b0;
    assign proc_6_data_PIPO_blk[18] = 1'b0;
    assign proc_6_start_FIFO_blk[18] = 1'b0;
    assign proc_6_TLF_FIFO_blk[18] = 1'b0;
    assign proc_6_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_6_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_6[18] = dl_detect_out ? proc_dep_vld_vec_6_reg[18] : (proc_6_data_FIFO_blk[18] | proc_6_data_PIPO_blk[18] | proc_6_start_FIFO_blk[18] | proc_6_TLF_FIFO_blk[18] | proc_6_input_sync_blk[18] | proc_6_output_sync_blk[18]);
    assign proc_6_data_FIFO_blk[19] = 1'b0;
    assign proc_6_data_PIPO_blk[19] = 1'b0;
    assign proc_6_start_FIFO_blk[19] = 1'b0;
    assign proc_6_TLF_FIFO_blk[19] = 1'b0;
    assign proc_6_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_6_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_6[19] = dl_detect_out ? proc_dep_vld_vec_6_reg[19] : (proc_6_data_FIFO_blk[19] | proc_6_data_PIPO_blk[19] | proc_6_start_FIFO_blk[19] | proc_6_TLF_FIFO_blk[19] | proc_6_input_sync_blk[19] | proc_6_output_sync_blk[19]);
    assign proc_6_data_FIFO_blk[20] = 1'b0;
    assign proc_6_data_PIPO_blk[20] = 1'b0;
    assign proc_6_start_FIFO_blk[20] = 1'b0;
    assign proc_6_TLF_FIFO_blk[20] = 1'b0;
    assign proc_6_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_6_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_6[20] = dl_detect_out ? proc_dep_vld_vec_6_reg[20] : (proc_6_data_FIFO_blk[20] | proc_6_data_PIPO_blk[20] | proc_6_start_FIFO_blk[20] | proc_6_TLF_FIFO_blk[20] | proc_6_input_sync_blk[20] | proc_6_output_sync_blk[20]);
    assign proc_6_data_FIFO_blk[21] = 1'b0;
    assign proc_6_data_PIPO_blk[21] = 1'b0;
    assign proc_6_start_FIFO_blk[21] = 1'b0;
    assign proc_6_TLF_FIFO_blk[21] = 1'b0;
    assign proc_6_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_6_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_6[21] = dl_detect_out ? proc_dep_vld_vec_6_reg[21] : (proc_6_data_FIFO_blk[21] | proc_6_data_PIPO_blk[21] | proc_6_start_FIFO_blk[21] | proc_6_TLF_FIFO_blk[21] | proc_6_input_sync_blk[21] | proc_6_output_sync_blk[21]);
    assign proc_6_data_FIFO_blk[22] = 1'b0;
    assign proc_6_data_PIPO_blk[22] = 1'b0;
    assign proc_6_start_FIFO_blk[22] = 1'b0;
    assign proc_6_TLF_FIFO_blk[22] = 1'b0;
    assign proc_6_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_6_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_6[22] = dl_detect_out ? proc_dep_vld_vec_6_reg[22] : (proc_6_data_FIFO_blk[22] | proc_6_data_PIPO_blk[22] | proc_6_start_FIFO_blk[22] | proc_6_TLF_FIFO_blk[22] | proc_6_input_sync_blk[22] | proc_6_output_sync_blk[22]);
    assign proc_6_data_FIFO_blk[23] = 1'b0;
    assign proc_6_data_PIPO_blk[23] = 1'b0;
    assign proc_6_start_FIFO_blk[23] = 1'b0;
    assign proc_6_TLF_FIFO_blk[23] = 1'b0;
    assign proc_6_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_6_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_6[23] = dl_detect_out ? proc_dep_vld_vec_6_reg[23] : (proc_6_data_FIFO_blk[23] | proc_6_data_PIPO_blk[23] | proc_6_start_FIFO_blk[23] | proc_6_TLF_FIFO_blk[23] | proc_6_input_sync_blk[23] | proc_6_output_sync_blk[23]);
    assign proc_6_data_FIFO_blk[24] = 1'b0;
    assign proc_6_data_PIPO_blk[24] = 1'b0;
    assign proc_6_start_FIFO_blk[24] = 1'b0;
    assign proc_6_TLF_FIFO_blk[24] = 1'b0;
    assign proc_6_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_6_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_6[24] = dl_detect_out ? proc_dep_vld_vec_6_reg[24] : (proc_6_data_FIFO_blk[24] | proc_6_data_PIPO_blk[24] | proc_6_start_FIFO_blk[24] | proc_6_TLF_FIFO_blk[24] | proc_6_input_sync_blk[24] | proc_6_output_sync_blk[24]);
    assign proc_6_data_FIFO_blk[25] = 1'b0;
    assign proc_6_data_PIPO_blk[25] = 1'b0;
    assign proc_6_start_FIFO_blk[25] = 1'b0;
    assign proc_6_TLF_FIFO_blk[25] = 1'b0;
    assign proc_6_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_6_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_6[25] = dl_detect_out ? proc_dep_vld_vec_6_reg[25] : (proc_6_data_FIFO_blk[25] | proc_6_data_PIPO_blk[25] | proc_6_start_FIFO_blk[25] | proc_6_TLF_FIFO_blk[25] | proc_6_input_sync_blk[25] | proc_6_output_sync_blk[25]);
    assign proc_6_data_FIFO_blk[26] = 1'b0;
    assign proc_6_data_PIPO_blk[26] = 1'b0;
    assign proc_6_start_FIFO_blk[26] = 1'b0;
    assign proc_6_TLF_FIFO_blk[26] = 1'b0;
    assign proc_6_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_6_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_6[26] = dl_detect_out ? proc_dep_vld_vec_6_reg[26] : (proc_6_data_FIFO_blk[26] | proc_6_data_PIPO_blk[26] | proc_6_start_FIFO_blk[26] | proc_6_TLF_FIFO_blk[26] | proc_6_input_sync_blk[26] | proc_6_output_sync_blk[26]);
    assign proc_6_data_FIFO_blk[27] = 1'b0;
    assign proc_6_data_PIPO_blk[27] = 1'b0;
    assign proc_6_start_FIFO_blk[27] = 1'b0;
    assign proc_6_TLF_FIFO_blk[27] = 1'b0;
    assign proc_6_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_6_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_6[27] = dl_detect_out ? proc_dep_vld_vec_6_reg[27] : (proc_6_data_FIFO_blk[27] | proc_6_data_PIPO_blk[27] | proc_6_start_FIFO_blk[27] | proc_6_TLF_FIFO_blk[27] | proc_6_input_sync_blk[27] | proc_6_output_sync_blk[27]);
    assign proc_6_data_FIFO_blk[28] = 1'b0;
    assign proc_6_data_PIPO_blk[28] = 1'b0;
    assign proc_6_start_FIFO_blk[28] = 1'b0;
    assign proc_6_TLF_FIFO_blk[28] = 1'b0;
    assign proc_6_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_6_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_6[28] = dl_detect_out ? proc_dep_vld_vec_6_reg[28] : (proc_6_data_FIFO_blk[28] | proc_6_data_PIPO_blk[28] | proc_6_start_FIFO_blk[28] | proc_6_TLF_FIFO_blk[28] | proc_6_input_sync_blk[28] | proc_6_output_sync_blk[28]);
    assign proc_6_data_FIFO_blk[29] = 1'b0;
    assign proc_6_data_PIPO_blk[29] = 1'b0;
    assign proc_6_start_FIFO_blk[29] = 1'b0;
    assign proc_6_TLF_FIFO_blk[29] = 1'b0;
    assign proc_6_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_6_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_6[29] = dl_detect_out ? proc_dep_vld_vec_6_reg[29] : (proc_6_data_FIFO_blk[29] | proc_6_data_PIPO_blk[29] | proc_6_start_FIFO_blk[29] | proc_6_TLF_FIFO_blk[29] | proc_6_input_sync_blk[29] | proc_6_output_sync_blk[29]);
    assign proc_6_data_FIFO_blk[30] = 1'b0;
    assign proc_6_data_PIPO_blk[30] = 1'b0;
    assign proc_6_start_FIFO_blk[30] = 1'b0;
    assign proc_6_TLF_FIFO_blk[30] = 1'b0;
    assign proc_6_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_6_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_6[30] = dl_detect_out ? proc_dep_vld_vec_6_reg[30] : (proc_6_data_FIFO_blk[30] | proc_6_data_PIPO_blk[30] | proc_6_start_FIFO_blk[30] | proc_6_TLF_FIFO_blk[30] | proc_6_input_sync_blk[30] | proc_6_output_sync_blk[30]);
    assign proc_6_data_FIFO_blk[31] = 1'b0;
    assign proc_6_data_PIPO_blk[31] = 1'b0;
    assign proc_6_start_FIFO_blk[31] = 1'b0;
    assign proc_6_TLF_FIFO_blk[31] = 1'b0;
    assign proc_6_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_6_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_6[31] = dl_detect_out ? proc_dep_vld_vec_6_reg[31] : (proc_6_data_FIFO_blk[31] | proc_6_data_PIPO_blk[31] | proc_6_start_FIFO_blk[31] | proc_6_TLF_FIFO_blk[31] | proc_6_input_sync_blk[31] | proc_6_output_sync_blk[31]);
    assign proc_6_data_FIFO_blk[32] = 1'b0;
    assign proc_6_data_PIPO_blk[32] = 1'b0;
    assign proc_6_start_FIFO_blk[32] = 1'b0;
    assign proc_6_TLF_FIFO_blk[32] = 1'b0;
    assign proc_6_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_6_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_6[32] = dl_detect_out ? proc_dep_vld_vec_6_reg[32] : (proc_6_data_FIFO_blk[32] | proc_6_data_PIPO_blk[32] | proc_6_start_FIFO_blk[32] | proc_6_TLF_FIFO_blk[32] | proc_6_input_sync_blk[32] | proc_6_output_sync_blk[32]);
    assign proc_6_data_FIFO_blk[33] = 1'b0;
    assign proc_6_data_PIPO_blk[33] = 1'b0;
    assign proc_6_start_FIFO_blk[33] = 1'b0;
    assign proc_6_TLF_FIFO_blk[33] = 1'b0;
    assign proc_6_input_sync_blk[33] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_6_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_6[33] = dl_detect_out ? proc_dep_vld_vec_6_reg[33] : (proc_6_data_FIFO_blk[33] | proc_6_data_PIPO_blk[33] | proc_6_start_FIFO_blk[33] | proc_6_TLF_FIFO_blk[33] | proc_6_input_sync_blk[33] | proc_6_output_sync_blk[33]);
    assign proc_6_data_FIFO_blk[34] = 1'b0;
    assign proc_6_data_PIPO_blk[34] = 1'b0;
    assign proc_6_start_FIFO_blk[34] = 1'b0;
    assign proc_6_TLF_FIFO_blk[34] = 1'b0;
    assign proc_6_input_sync_blk[34] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_6_output_sync_blk[34] = 1'b0;
    assign proc_dep_vld_vec_6[34] = dl_detect_out ? proc_dep_vld_vec_6_reg[34] : (proc_6_data_FIFO_blk[34] | proc_6_data_PIPO_blk[34] | proc_6_start_FIFO_blk[34] | proc_6_TLF_FIFO_blk[34] | proc_6_input_sync_blk[34] | proc_6_output_sync_blk[34]);
    assign proc_6_data_FIFO_blk[35] = 1'b0;
    assign proc_6_data_PIPO_blk[35] = 1'b0;
    assign proc_6_start_FIFO_blk[35] = 1'b0;
    assign proc_6_TLF_FIFO_blk[35] = 1'b0;
    assign proc_6_input_sync_blk[35] = 1'b0 | (ap_sync_ProcessingElement_1_U0_ap_ready & ProcessingElement_1_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_6_output_sync_blk[35] = 1'b0;
    assign proc_dep_vld_vec_6[35] = dl_detect_out ? proc_dep_vld_vec_6_reg[35] : (proc_6_data_FIFO_blk[35] | proc_6_data_PIPO_blk[35] | proc_6_start_FIFO_blk[35] | proc_6_TLF_FIFO_blk[35] | proc_6_input_sync_blk[35] | proc_6_output_sync_blk[35]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_6_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_6_reg <= proc_dep_vld_vec_6;
        end
    end
    assign in_chan_dep_vld_vec_6[0] = dep_chan_vld_0_6;
    assign in_chan_dep_data_vec_6[39 : 0] = dep_chan_data_0_6;
    assign token_in_vec_6[0] = token_0_6;
    assign in_chan_dep_vld_vec_6[1] = dep_chan_vld_1_6;
    assign in_chan_dep_data_vec_6[79 : 40] = dep_chan_data_1_6;
    assign token_in_vec_6[1] = token_1_6;
    assign in_chan_dep_vld_vec_6[2] = dep_chan_vld_2_6;
    assign in_chan_dep_data_vec_6[119 : 80] = dep_chan_data_2_6;
    assign token_in_vec_6[2] = token_2_6;
    assign in_chan_dep_vld_vec_6[3] = dep_chan_vld_3_6;
    assign in_chan_dep_data_vec_6[159 : 120] = dep_chan_data_3_6;
    assign token_in_vec_6[3] = token_3_6;
    assign in_chan_dep_vld_vec_6[4] = dep_chan_vld_5_6;
    assign in_chan_dep_data_vec_6[199 : 160] = dep_chan_data_5_6;
    assign token_in_vec_6[4] = token_5_6;
    assign in_chan_dep_vld_vec_6[5] = dep_chan_vld_7_6;
    assign in_chan_dep_data_vec_6[239 : 200] = dep_chan_data_7_6;
    assign token_in_vec_6[5] = token_7_6;
    assign in_chan_dep_vld_vec_6[6] = dep_chan_vld_8_6;
    assign in_chan_dep_data_vec_6[279 : 240] = dep_chan_data_8_6;
    assign token_in_vec_6[6] = token_8_6;
    assign in_chan_dep_vld_vec_6[7] = dep_chan_vld_9_6;
    assign in_chan_dep_data_vec_6[319 : 280] = dep_chan_data_9_6;
    assign token_in_vec_6[7] = token_9_6;
    assign in_chan_dep_vld_vec_6[8] = dep_chan_vld_10_6;
    assign in_chan_dep_data_vec_6[359 : 320] = dep_chan_data_10_6;
    assign token_in_vec_6[8] = token_10_6;
    assign in_chan_dep_vld_vec_6[9] = dep_chan_vld_11_6;
    assign in_chan_dep_data_vec_6[399 : 360] = dep_chan_data_11_6;
    assign token_in_vec_6[9] = token_11_6;
    assign in_chan_dep_vld_vec_6[10] = dep_chan_vld_12_6;
    assign in_chan_dep_data_vec_6[439 : 400] = dep_chan_data_12_6;
    assign token_in_vec_6[10] = token_12_6;
    assign in_chan_dep_vld_vec_6[11] = dep_chan_vld_13_6;
    assign in_chan_dep_data_vec_6[479 : 440] = dep_chan_data_13_6;
    assign token_in_vec_6[11] = token_13_6;
    assign in_chan_dep_vld_vec_6[12] = dep_chan_vld_14_6;
    assign in_chan_dep_data_vec_6[519 : 480] = dep_chan_data_14_6;
    assign token_in_vec_6[12] = token_14_6;
    assign in_chan_dep_vld_vec_6[13] = dep_chan_vld_15_6;
    assign in_chan_dep_data_vec_6[559 : 520] = dep_chan_data_15_6;
    assign token_in_vec_6[13] = token_15_6;
    assign in_chan_dep_vld_vec_6[14] = dep_chan_vld_16_6;
    assign in_chan_dep_data_vec_6[599 : 560] = dep_chan_data_16_6;
    assign token_in_vec_6[14] = token_16_6;
    assign in_chan_dep_vld_vec_6[15] = dep_chan_vld_17_6;
    assign in_chan_dep_data_vec_6[639 : 600] = dep_chan_data_17_6;
    assign token_in_vec_6[15] = token_17_6;
    assign in_chan_dep_vld_vec_6[16] = dep_chan_vld_18_6;
    assign in_chan_dep_data_vec_6[679 : 640] = dep_chan_data_18_6;
    assign token_in_vec_6[16] = token_18_6;
    assign in_chan_dep_vld_vec_6[17] = dep_chan_vld_19_6;
    assign in_chan_dep_data_vec_6[719 : 680] = dep_chan_data_19_6;
    assign token_in_vec_6[17] = token_19_6;
    assign in_chan_dep_vld_vec_6[18] = dep_chan_vld_20_6;
    assign in_chan_dep_data_vec_6[759 : 720] = dep_chan_data_20_6;
    assign token_in_vec_6[18] = token_20_6;
    assign in_chan_dep_vld_vec_6[19] = dep_chan_vld_21_6;
    assign in_chan_dep_data_vec_6[799 : 760] = dep_chan_data_21_6;
    assign token_in_vec_6[19] = token_21_6;
    assign in_chan_dep_vld_vec_6[20] = dep_chan_vld_22_6;
    assign in_chan_dep_data_vec_6[839 : 800] = dep_chan_data_22_6;
    assign token_in_vec_6[20] = token_22_6;
    assign in_chan_dep_vld_vec_6[21] = dep_chan_vld_23_6;
    assign in_chan_dep_data_vec_6[879 : 840] = dep_chan_data_23_6;
    assign token_in_vec_6[21] = token_23_6;
    assign in_chan_dep_vld_vec_6[22] = dep_chan_vld_24_6;
    assign in_chan_dep_data_vec_6[919 : 880] = dep_chan_data_24_6;
    assign token_in_vec_6[22] = token_24_6;
    assign in_chan_dep_vld_vec_6[23] = dep_chan_vld_25_6;
    assign in_chan_dep_data_vec_6[959 : 920] = dep_chan_data_25_6;
    assign token_in_vec_6[23] = token_25_6;
    assign in_chan_dep_vld_vec_6[24] = dep_chan_vld_26_6;
    assign in_chan_dep_data_vec_6[999 : 960] = dep_chan_data_26_6;
    assign token_in_vec_6[24] = token_26_6;
    assign in_chan_dep_vld_vec_6[25] = dep_chan_vld_27_6;
    assign in_chan_dep_data_vec_6[1039 : 1000] = dep_chan_data_27_6;
    assign token_in_vec_6[25] = token_27_6;
    assign in_chan_dep_vld_vec_6[26] = dep_chan_vld_28_6;
    assign in_chan_dep_data_vec_6[1079 : 1040] = dep_chan_data_28_6;
    assign token_in_vec_6[26] = token_28_6;
    assign in_chan_dep_vld_vec_6[27] = dep_chan_vld_29_6;
    assign in_chan_dep_data_vec_6[1119 : 1080] = dep_chan_data_29_6;
    assign token_in_vec_6[27] = token_29_6;
    assign in_chan_dep_vld_vec_6[28] = dep_chan_vld_30_6;
    assign in_chan_dep_data_vec_6[1159 : 1120] = dep_chan_data_30_6;
    assign token_in_vec_6[28] = token_30_6;
    assign in_chan_dep_vld_vec_6[29] = dep_chan_vld_31_6;
    assign in_chan_dep_data_vec_6[1199 : 1160] = dep_chan_data_31_6;
    assign token_in_vec_6[29] = token_31_6;
    assign in_chan_dep_vld_vec_6[30] = dep_chan_vld_32_6;
    assign in_chan_dep_data_vec_6[1239 : 1200] = dep_chan_data_32_6;
    assign token_in_vec_6[30] = token_32_6;
    assign in_chan_dep_vld_vec_6[31] = dep_chan_vld_33_6;
    assign in_chan_dep_data_vec_6[1279 : 1240] = dep_chan_data_33_6;
    assign token_in_vec_6[31] = token_33_6;
    assign in_chan_dep_vld_vec_6[32] = dep_chan_vld_34_6;
    assign in_chan_dep_data_vec_6[1319 : 1280] = dep_chan_data_34_6;
    assign token_in_vec_6[32] = token_34_6;
    assign in_chan_dep_vld_vec_6[33] = dep_chan_vld_35_6;
    assign in_chan_dep_data_vec_6[1359 : 1320] = dep_chan_data_35_6;
    assign token_in_vec_6[33] = token_35_6;
    assign in_chan_dep_vld_vec_6[34] = dep_chan_vld_36_6;
    assign in_chan_dep_data_vec_6[1399 : 1360] = dep_chan_data_36_6;
    assign token_in_vec_6[34] = token_36_6;
    assign in_chan_dep_vld_vec_6[35] = dep_chan_vld_38_6;
    assign in_chan_dep_data_vec_6[1439 : 1400] = dep_chan_data_38_6;
    assign token_in_vec_6[35] = token_38_6;
    assign dep_chan_vld_6_2 = out_chan_dep_vld_vec_6[0];
    assign dep_chan_data_6_2 = out_chan_dep_data_6;
    assign token_6_2 = token_out_vec_6[0];
    assign dep_chan_vld_6_7 = out_chan_dep_vld_vec_6[1];
    assign dep_chan_data_6_7 = out_chan_dep_data_6;
    assign token_6_7 = token_out_vec_6[1];
    assign dep_chan_vld_6_5 = out_chan_dep_vld_vec_6[2];
    assign dep_chan_data_6_5 = out_chan_dep_data_6;
    assign token_6_5 = token_out_vec_6[2];
    assign dep_chan_vld_6_38 = out_chan_dep_vld_vec_6[3];
    assign dep_chan_data_6_38 = out_chan_dep_data_6;
    assign token_6_38 = token_out_vec_6[3];
    assign dep_chan_vld_6_0 = out_chan_dep_vld_vec_6[4];
    assign dep_chan_data_6_0 = out_chan_dep_data_6;
    assign token_6_0 = token_out_vec_6[4];
    assign dep_chan_vld_6_1 = out_chan_dep_vld_vec_6[5];
    assign dep_chan_data_6_1 = out_chan_dep_data_6;
    assign token_6_1 = token_out_vec_6[5];
    assign dep_chan_vld_6_3 = out_chan_dep_vld_vec_6[6];
    assign dep_chan_data_6_3 = out_chan_dep_data_6;
    assign token_6_3 = token_out_vec_6[6];
    assign dep_chan_vld_6_8 = out_chan_dep_vld_vec_6[7];
    assign dep_chan_data_6_8 = out_chan_dep_data_6;
    assign token_6_8 = token_out_vec_6[7];
    assign dep_chan_vld_6_9 = out_chan_dep_vld_vec_6[8];
    assign dep_chan_data_6_9 = out_chan_dep_data_6;
    assign token_6_9 = token_out_vec_6[8];
    assign dep_chan_vld_6_10 = out_chan_dep_vld_vec_6[9];
    assign dep_chan_data_6_10 = out_chan_dep_data_6;
    assign token_6_10 = token_out_vec_6[9];
    assign dep_chan_vld_6_11 = out_chan_dep_vld_vec_6[10];
    assign dep_chan_data_6_11 = out_chan_dep_data_6;
    assign token_6_11 = token_out_vec_6[10];
    assign dep_chan_vld_6_12 = out_chan_dep_vld_vec_6[11];
    assign dep_chan_data_6_12 = out_chan_dep_data_6;
    assign token_6_12 = token_out_vec_6[11];
    assign dep_chan_vld_6_13 = out_chan_dep_vld_vec_6[12];
    assign dep_chan_data_6_13 = out_chan_dep_data_6;
    assign token_6_13 = token_out_vec_6[12];
    assign dep_chan_vld_6_14 = out_chan_dep_vld_vec_6[13];
    assign dep_chan_data_6_14 = out_chan_dep_data_6;
    assign token_6_14 = token_out_vec_6[13];
    assign dep_chan_vld_6_15 = out_chan_dep_vld_vec_6[14];
    assign dep_chan_data_6_15 = out_chan_dep_data_6;
    assign token_6_15 = token_out_vec_6[14];
    assign dep_chan_vld_6_16 = out_chan_dep_vld_vec_6[15];
    assign dep_chan_data_6_16 = out_chan_dep_data_6;
    assign token_6_16 = token_out_vec_6[15];
    assign dep_chan_vld_6_17 = out_chan_dep_vld_vec_6[16];
    assign dep_chan_data_6_17 = out_chan_dep_data_6;
    assign token_6_17 = token_out_vec_6[16];
    assign dep_chan_vld_6_18 = out_chan_dep_vld_vec_6[17];
    assign dep_chan_data_6_18 = out_chan_dep_data_6;
    assign token_6_18 = token_out_vec_6[17];
    assign dep_chan_vld_6_19 = out_chan_dep_vld_vec_6[18];
    assign dep_chan_data_6_19 = out_chan_dep_data_6;
    assign token_6_19 = token_out_vec_6[18];
    assign dep_chan_vld_6_20 = out_chan_dep_vld_vec_6[19];
    assign dep_chan_data_6_20 = out_chan_dep_data_6;
    assign token_6_20 = token_out_vec_6[19];
    assign dep_chan_vld_6_21 = out_chan_dep_vld_vec_6[20];
    assign dep_chan_data_6_21 = out_chan_dep_data_6;
    assign token_6_21 = token_out_vec_6[20];
    assign dep_chan_vld_6_22 = out_chan_dep_vld_vec_6[21];
    assign dep_chan_data_6_22 = out_chan_dep_data_6;
    assign token_6_22 = token_out_vec_6[21];
    assign dep_chan_vld_6_23 = out_chan_dep_vld_vec_6[22];
    assign dep_chan_data_6_23 = out_chan_dep_data_6;
    assign token_6_23 = token_out_vec_6[22];
    assign dep_chan_vld_6_24 = out_chan_dep_vld_vec_6[23];
    assign dep_chan_data_6_24 = out_chan_dep_data_6;
    assign token_6_24 = token_out_vec_6[23];
    assign dep_chan_vld_6_25 = out_chan_dep_vld_vec_6[24];
    assign dep_chan_data_6_25 = out_chan_dep_data_6;
    assign token_6_25 = token_out_vec_6[24];
    assign dep_chan_vld_6_26 = out_chan_dep_vld_vec_6[25];
    assign dep_chan_data_6_26 = out_chan_dep_data_6;
    assign token_6_26 = token_out_vec_6[25];
    assign dep_chan_vld_6_27 = out_chan_dep_vld_vec_6[26];
    assign dep_chan_data_6_27 = out_chan_dep_data_6;
    assign token_6_27 = token_out_vec_6[26];
    assign dep_chan_vld_6_28 = out_chan_dep_vld_vec_6[27];
    assign dep_chan_data_6_28 = out_chan_dep_data_6;
    assign token_6_28 = token_out_vec_6[27];
    assign dep_chan_vld_6_29 = out_chan_dep_vld_vec_6[28];
    assign dep_chan_data_6_29 = out_chan_dep_data_6;
    assign token_6_29 = token_out_vec_6[28];
    assign dep_chan_vld_6_30 = out_chan_dep_vld_vec_6[29];
    assign dep_chan_data_6_30 = out_chan_dep_data_6;
    assign token_6_30 = token_out_vec_6[29];
    assign dep_chan_vld_6_31 = out_chan_dep_vld_vec_6[30];
    assign dep_chan_data_6_31 = out_chan_dep_data_6;
    assign token_6_31 = token_out_vec_6[30];
    assign dep_chan_vld_6_32 = out_chan_dep_vld_vec_6[31];
    assign dep_chan_data_6_32 = out_chan_dep_data_6;
    assign token_6_32 = token_out_vec_6[31];
    assign dep_chan_vld_6_33 = out_chan_dep_vld_vec_6[32];
    assign dep_chan_data_6_33 = out_chan_dep_data_6;
    assign token_6_33 = token_out_vec_6[32];
    assign dep_chan_vld_6_34 = out_chan_dep_vld_vec_6[33];
    assign dep_chan_data_6_34 = out_chan_dep_data_6;
    assign token_6_34 = token_out_vec_6[33];
    assign dep_chan_vld_6_35 = out_chan_dep_vld_vec_6[34];
    assign dep_chan_data_6_35 = out_chan_dep_data_6;
    assign token_6_35 = token_out_vec_6[34];
    assign dep_chan_vld_6_36 = out_chan_dep_vld_vec_6[35];
    assign dep_chan_data_6_36 = out_chan_dep_data_6;
    assign token_6_36 = token_out_vec_6[35];

    // Process: ProcessingElement_2_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 7, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_7 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_7),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_7),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_7),
        .token_in_vec(token_in_vec_7),
        .dl_detect_in(dl_detect_out),
        .origin(origin[7]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_7),
        .out_chan_dep_data(out_chan_dep_data_7),
        .token_out_vec(token_out_vec_7),
        .dl_detect_out(dl_in_vec[7]));

    assign proc_7_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_1_blk_n) | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_1_blk_n) | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_WriteC_Flattened_fu_179.cPipes_1_blk_n);
    assign proc_7_data_PIPO_blk[0] = 1'b0;
    assign proc_7_start_FIFO_blk[0] = 1'b0;
    assign proc_7_TLF_FIFO_blk[0] = 1'b0;
    assign proc_7_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_7_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_7[0] = dl_detect_out ? proc_dep_vld_vec_7_reg[0] : (proc_7_data_FIFO_blk[0] | proc_7_data_PIPO_blk[0] | proc_7_start_FIFO_blk[0] | proc_7_TLF_FIFO_blk[0] | proc_7_input_sync_blk[0] | proc_7_output_sync_blk[0]);
    assign proc_7_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_2_blk_n) | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_2_blk_n) | (~ProcessingElement_2_U0.grp_ProcessingElement_2_Pipeline_WriteC_Flattened_fu_179.cPipes_2_blk_n);
    assign proc_7_data_PIPO_blk[1] = 1'b0;
    assign proc_7_start_FIFO_blk[1] = 1'b0;
    assign proc_7_TLF_FIFO_blk[1] = 1'b0;
    assign proc_7_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_7_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_7[1] = dl_detect_out ? proc_dep_vld_vec_7_reg[1] : (proc_7_data_FIFO_blk[1] | proc_7_data_PIPO_blk[1] | proc_7_start_FIFO_blk[1] | proc_7_TLF_FIFO_blk[1] | proc_7_input_sync_blk[1] | proc_7_output_sync_blk[1]);
    assign proc_7_data_FIFO_blk[2] = 1'b0;
    assign proc_7_data_PIPO_blk[2] = 1'b0;
    assign proc_7_start_FIFO_blk[2] = 1'b0;
    assign proc_7_TLF_FIFO_blk[2] = 1'b0;
    assign proc_7_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_7_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_7[2] = dl_detect_out ? proc_dep_vld_vec_7_reg[2] : (proc_7_data_FIFO_blk[2] | proc_7_data_PIPO_blk[2] | proc_7_start_FIFO_blk[2] | proc_7_TLF_FIFO_blk[2] | proc_7_input_sync_blk[2] | proc_7_output_sync_blk[2]);
    assign proc_7_data_FIFO_blk[3] = 1'b0;
    assign proc_7_data_PIPO_blk[3] = 1'b0;
    assign proc_7_start_FIFO_blk[3] = 1'b0;
    assign proc_7_TLF_FIFO_blk[3] = 1'b0;
    assign proc_7_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_7_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_7[3] = dl_detect_out ? proc_dep_vld_vec_7_reg[3] : (proc_7_data_FIFO_blk[3] | proc_7_data_PIPO_blk[3] | proc_7_start_FIFO_blk[3] | proc_7_TLF_FIFO_blk[3] | proc_7_input_sync_blk[3] | proc_7_output_sync_blk[3]);
    assign proc_7_data_FIFO_blk[4] = 1'b0;
    assign proc_7_data_PIPO_blk[4] = 1'b0;
    assign proc_7_start_FIFO_blk[4] = 1'b0;
    assign proc_7_TLF_FIFO_blk[4] = 1'b0;
    assign proc_7_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_7_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_7[4] = dl_detect_out ? proc_dep_vld_vec_7_reg[4] : (proc_7_data_FIFO_blk[4] | proc_7_data_PIPO_blk[4] | proc_7_start_FIFO_blk[4] | proc_7_TLF_FIFO_blk[4] | proc_7_input_sync_blk[4] | proc_7_output_sync_blk[4]);
    assign proc_7_data_FIFO_blk[5] = 1'b0;
    assign proc_7_data_PIPO_blk[5] = 1'b0;
    assign proc_7_start_FIFO_blk[5] = 1'b0;
    assign proc_7_TLF_FIFO_blk[5] = 1'b0;
    assign proc_7_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_7_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_7[5] = dl_detect_out ? proc_dep_vld_vec_7_reg[5] : (proc_7_data_FIFO_blk[5] | proc_7_data_PIPO_blk[5] | proc_7_start_FIFO_blk[5] | proc_7_TLF_FIFO_blk[5] | proc_7_input_sync_blk[5] | proc_7_output_sync_blk[5]);
    assign proc_7_data_FIFO_blk[6] = 1'b0;
    assign proc_7_data_PIPO_blk[6] = 1'b0;
    assign proc_7_start_FIFO_blk[6] = 1'b0;
    assign proc_7_TLF_FIFO_blk[6] = 1'b0;
    assign proc_7_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_7_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_7[6] = dl_detect_out ? proc_dep_vld_vec_7_reg[6] : (proc_7_data_FIFO_blk[6] | proc_7_data_PIPO_blk[6] | proc_7_start_FIFO_blk[6] | proc_7_TLF_FIFO_blk[6] | proc_7_input_sync_blk[6] | proc_7_output_sync_blk[6]);
    assign proc_7_data_FIFO_blk[7] = 1'b0;
    assign proc_7_data_PIPO_blk[7] = 1'b0;
    assign proc_7_start_FIFO_blk[7] = 1'b0;
    assign proc_7_TLF_FIFO_blk[7] = 1'b0;
    assign proc_7_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_7_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_7[7] = dl_detect_out ? proc_dep_vld_vec_7_reg[7] : (proc_7_data_FIFO_blk[7] | proc_7_data_PIPO_blk[7] | proc_7_start_FIFO_blk[7] | proc_7_TLF_FIFO_blk[7] | proc_7_input_sync_blk[7] | proc_7_output_sync_blk[7]);
    assign proc_7_data_FIFO_blk[8] = 1'b0;
    assign proc_7_data_PIPO_blk[8] = 1'b0;
    assign proc_7_start_FIFO_blk[8] = 1'b0;
    assign proc_7_TLF_FIFO_blk[8] = 1'b0;
    assign proc_7_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_7_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_7[8] = dl_detect_out ? proc_dep_vld_vec_7_reg[8] : (proc_7_data_FIFO_blk[8] | proc_7_data_PIPO_blk[8] | proc_7_start_FIFO_blk[8] | proc_7_TLF_FIFO_blk[8] | proc_7_input_sync_blk[8] | proc_7_output_sync_blk[8]);
    assign proc_7_data_FIFO_blk[9] = 1'b0;
    assign proc_7_data_PIPO_blk[9] = 1'b0;
    assign proc_7_start_FIFO_blk[9] = 1'b0;
    assign proc_7_TLF_FIFO_blk[9] = 1'b0;
    assign proc_7_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_7_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_7[9] = dl_detect_out ? proc_dep_vld_vec_7_reg[9] : (proc_7_data_FIFO_blk[9] | proc_7_data_PIPO_blk[9] | proc_7_start_FIFO_blk[9] | proc_7_TLF_FIFO_blk[9] | proc_7_input_sync_blk[9] | proc_7_output_sync_blk[9]);
    assign proc_7_data_FIFO_blk[10] = 1'b0;
    assign proc_7_data_PIPO_blk[10] = 1'b0;
    assign proc_7_start_FIFO_blk[10] = 1'b0;
    assign proc_7_TLF_FIFO_blk[10] = 1'b0;
    assign proc_7_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_7_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_7[10] = dl_detect_out ? proc_dep_vld_vec_7_reg[10] : (proc_7_data_FIFO_blk[10] | proc_7_data_PIPO_blk[10] | proc_7_start_FIFO_blk[10] | proc_7_TLF_FIFO_blk[10] | proc_7_input_sync_blk[10] | proc_7_output_sync_blk[10]);
    assign proc_7_data_FIFO_blk[11] = 1'b0;
    assign proc_7_data_PIPO_blk[11] = 1'b0;
    assign proc_7_start_FIFO_blk[11] = 1'b0;
    assign proc_7_TLF_FIFO_blk[11] = 1'b0;
    assign proc_7_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_7_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_7[11] = dl_detect_out ? proc_dep_vld_vec_7_reg[11] : (proc_7_data_FIFO_blk[11] | proc_7_data_PIPO_blk[11] | proc_7_start_FIFO_blk[11] | proc_7_TLF_FIFO_blk[11] | proc_7_input_sync_blk[11] | proc_7_output_sync_blk[11]);
    assign proc_7_data_FIFO_blk[12] = 1'b0;
    assign proc_7_data_PIPO_blk[12] = 1'b0;
    assign proc_7_start_FIFO_blk[12] = 1'b0;
    assign proc_7_TLF_FIFO_blk[12] = 1'b0;
    assign proc_7_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_7_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_7[12] = dl_detect_out ? proc_dep_vld_vec_7_reg[12] : (proc_7_data_FIFO_blk[12] | proc_7_data_PIPO_blk[12] | proc_7_start_FIFO_blk[12] | proc_7_TLF_FIFO_blk[12] | proc_7_input_sync_blk[12] | proc_7_output_sync_blk[12]);
    assign proc_7_data_FIFO_blk[13] = 1'b0;
    assign proc_7_data_PIPO_blk[13] = 1'b0;
    assign proc_7_start_FIFO_blk[13] = 1'b0;
    assign proc_7_TLF_FIFO_blk[13] = 1'b0;
    assign proc_7_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_7_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_7[13] = dl_detect_out ? proc_dep_vld_vec_7_reg[13] : (proc_7_data_FIFO_blk[13] | proc_7_data_PIPO_blk[13] | proc_7_start_FIFO_blk[13] | proc_7_TLF_FIFO_blk[13] | proc_7_input_sync_blk[13] | proc_7_output_sync_blk[13]);
    assign proc_7_data_FIFO_blk[14] = 1'b0;
    assign proc_7_data_PIPO_blk[14] = 1'b0;
    assign proc_7_start_FIFO_blk[14] = 1'b0;
    assign proc_7_TLF_FIFO_blk[14] = 1'b0;
    assign proc_7_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_7_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_7[14] = dl_detect_out ? proc_dep_vld_vec_7_reg[14] : (proc_7_data_FIFO_blk[14] | proc_7_data_PIPO_blk[14] | proc_7_start_FIFO_blk[14] | proc_7_TLF_FIFO_blk[14] | proc_7_input_sync_blk[14] | proc_7_output_sync_blk[14]);
    assign proc_7_data_FIFO_blk[15] = 1'b0;
    assign proc_7_data_PIPO_blk[15] = 1'b0;
    assign proc_7_start_FIFO_blk[15] = 1'b0;
    assign proc_7_TLF_FIFO_blk[15] = 1'b0;
    assign proc_7_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_7_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_7[15] = dl_detect_out ? proc_dep_vld_vec_7_reg[15] : (proc_7_data_FIFO_blk[15] | proc_7_data_PIPO_blk[15] | proc_7_start_FIFO_blk[15] | proc_7_TLF_FIFO_blk[15] | proc_7_input_sync_blk[15] | proc_7_output_sync_blk[15]);
    assign proc_7_data_FIFO_blk[16] = 1'b0;
    assign proc_7_data_PIPO_blk[16] = 1'b0;
    assign proc_7_start_FIFO_blk[16] = 1'b0;
    assign proc_7_TLF_FIFO_blk[16] = 1'b0;
    assign proc_7_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_7_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_7[16] = dl_detect_out ? proc_dep_vld_vec_7_reg[16] : (proc_7_data_FIFO_blk[16] | proc_7_data_PIPO_blk[16] | proc_7_start_FIFO_blk[16] | proc_7_TLF_FIFO_blk[16] | proc_7_input_sync_blk[16] | proc_7_output_sync_blk[16]);
    assign proc_7_data_FIFO_blk[17] = 1'b0;
    assign proc_7_data_PIPO_blk[17] = 1'b0;
    assign proc_7_start_FIFO_blk[17] = 1'b0;
    assign proc_7_TLF_FIFO_blk[17] = 1'b0;
    assign proc_7_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_7_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_7[17] = dl_detect_out ? proc_dep_vld_vec_7_reg[17] : (proc_7_data_FIFO_blk[17] | proc_7_data_PIPO_blk[17] | proc_7_start_FIFO_blk[17] | proc_7_TLF_FIFO_blk[17] | proc_7_input_sync_blk[17] | proc_7_output_sync_blk[17]);
    assign proc_7_data_FIFO_blk[18] = 1'b0;
    assign proc_7_data_PIPO_blk[18] = 1'b0;
    assign proc_7_start_FIFO_blk[18] = 1'b0;
    assign proc_7_TLF_FIFO_blk[18] = 1'b0;
    assign proc_7_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_7_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_7[18] = dl_detect_out ? proc_dep_vld_vec_7_reg[18] : (proc_7_data_FIFO_blk[18] | proc_7_data_PIPO_blk[18] | proc_7_start_FIFO_blk[18] | proc_7_TLF_FIFO_blk[18] | proc_7_input_sync_blk[18] | proc_7_output_sync_blk[18]);
    assign proc_7_data_FIFO_blk[19] = 1'b0;
    assign proc_7_data_PIPO_blk[19] = 1'b0;
    assign proc_7_start_FIFO_blk[19] = 1'b0;
    assign proc_7_TLF_FIFO_blk[19] = 1'b0;
    assign proc_7_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_7_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_7[19] = dl_detect_out ? proc_dep_vld_vec_7_reg[19] : (proc_7_data_FIFO_blk[19] | proc_7_data_PIPO_blk[19] | proc_7_start_FIFO_blk[19] | proc_7_TLF_FIFO_blk[19] | proc_7_input_sync_blk[19] | proc_7_output_sync_blk[19]);
    assign proc_7_data_FIFO_blk[20] = 1'b0;
    assign proc_7_data_PIPO_blk[20] = 1'b0;
    assign proc_7_start_FIFO_blk[20] = 1'b0;
    assign proc_7_TLF_FIFO_blk[20] = 1'b0;
    assign proc_7_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_7_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_7[20] = dl_detect_out ? proc_dep_vld_vec_7_reg[20] : (proc_7_data_FIFO_blk[20] | proc_7_data_PIPO_blk[20] | proc_7_start_FIFO_blk[20] | proc_7_TLF_FIFO_blk[20] | proc_7_input_sync_blk[20] | proc_7_output_sync_blk[20]);
    assign proc_7_data_FIFO_blk[21] = 1'b0;
    assign proc_7_data_PIPO_blk[21] = 1'b0;
    assign proc_7_start_FIFO_blk[21] = 1'b0;
    assign proc_7_TLF_FIFO_blk[21] = 1'b0;
    assign proc_7_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_7_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_7[21] = dl_detect_out ? proc_dep_vld_vec_7_reg[21] : (proc_7_data_FIFO_blk[21] | proc_7_data_PIPO_blk[21] | proc_7_start_FIFO_blk[21] | proc_7_TLF_FIFO_blk[21] | proc_7_input_sync_blk[21] | proc_7_output_sync_blk[21]);
    assign proc_7_data_FIFO_blk[22] = 1'b0;
    assign proc_7_data_PIPO_blk[22] = 1'b0;
    assign proc_7_start_FIFO_blk[22] = 1'b0;
    assign proc_7_TLF_FIFO_blk[22] = 1'b0;
    assign proc_7_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_7_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_7[22] = dl_detect_out ? proc_dep_vld_vec_7_reg[22] : (proc_7_data_FIFO_blk[22] | proc_7_data_PIPO_blk[22] | proc_7_start_FIFO_blk[22] | proc_7_TLF_FIFO_blk[22] | proc_7_input_sync_blk[22] | proc_7_output_sync_blk[22]);
    assign proc_7_data_FIFO_blk[23] = 1'b0;
    assign proc_7_data_PIPO_blk[23] = 1'b0;
    assign proc_7_start_FIFO_blk[23] = 1'b0;
    assign proc_7_TLF_FIFO_blk[23] = 1'b0;
    assign proc_7_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_7_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_7[23] = dl_detect_out ? proc_dep_vld_vec_7_reg[23] : (proc_7_data_FIFO_blk[23] | proc_7_data_PIPO_blk[23] | proc_7_start_FIFO_blk[23] | proc_7_TLF_FIFO_blk[23] | proc_7_input_sync_blk[23] | proc_7_output_sync_blk[23]);
    assign proc_7_data_FIFO_blk[24] = 1'b0;
    assign proc_7_data_PIPO_blk[24] = 1'b0;
    assign proc_7_start_FIFO_blk[24] = 1'b0;
    assign proc_7_TLF_FIFO_blk[24] = 1'b0;
    assign proc_7_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_7_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_7[24] = dl_detect_out ? proc_dep_vld_vec_7_reg[24] : (proc_7_data_FIFO_blk[24] | proc_7_data_PIPO_blk[24] | proc_7_start_FIFO_blk[24] | proc_7_TLF_FIFO_blk[24] | proc_7_input_sync_blk[24] | proc_7_output_sync_blk[24]);
    assign proc_7_data_FIFO_blk[25] = 1'b0;
    assign proc_7_data_PIPO_blk[25] = 1'b0;
    assign proc_7_start_FIFO_blk[25] = 1'b0;
    assign proc_7_TLF_FIFO_blk[25] = 1'b0;
    assign proc_7_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_7_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_7[25] = dl_detect_out ? proc_dep_vld_vec_7_reg[25] : (proc_7_data_FIFO_blk[25] | proc_7_data_PIPO_blk[25] | proc_7_start_FIFO_blk[25] | proc_7_TLF_FIFO_blk[25] | proc_7_input_sync_blk[25] | proc_7_output_sync_blk[25]);
    assign proc_7_data_FIFO_blk[26] = 1'b0;
    assign proc_7_data_PIPO_blk[26] = 1'b0;
    assign proc_7_start_FIFO_blk[26] = 1'b0;
    assign proc_7_TLF_FIFO_blk[26] = 1'b0;
    assign proc_7_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_7_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_7[26] = dl_detect_out ? proc_dep_vld_vec_7_reg[26] : (proc_7_data_FIFO_blk[26] | proc_7_data_PIPO_blk[26] | proc_7_start_FIFO_blk[26] | proc_7_TLF_FIFO_blk[26] | proc_7_input_sync_blk[26] | proc_7_output_sync_blk[26]);
    assign proc_7_data_FIFO_blk[27] = 1'b0;
    assign proc_7_data_PIPO_blk[27] = 1'b0;
    assign proc_7_start_FIFO_blk[27] = 1'b0;
    assign proc_7_TLF_FIFO_blk[27] = 1'b0;
    assign proc_7_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_7_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_7[27] = dl_detect_out ? proc_dep_vld_vec_7_reg[27] : (proc_7_data_FIFO_blk[27] | proc_7_data_PIPO_blk[27] | proc_7_start_FIFO_blk[27] | proc_7_TLF_FIFO_blk[27] | proc_7_input_sync_blk[27] | proc_7_output_sync_blk[27]);
    assign proc_7_data_FIFO_blk[28] = 1'b0;
    assign proc_7_data_PIPO_blk[28] = 1'b0;
    assign proc_7_start_FIFO_blk[28] = 1'b0;
    assign proc_7_TLF_FIFO_blk[28] = 1'b0;
    assign proc_7_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_7_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_7[28] = dl_detect_out ? proc_dep_vld_vec_7_reg[28] : (proc_7_data_FIFO_blk[28] | proc_7_data_PIPO_blk[28] | proc_7_start_FIFO_blk[28] | proc_7_TLF_FIFO_blk[28] | proc_7_input_sync_blk[28] | proc_7_output_sync_blk[28]);
    assign proc_7_data_FIFO_blk[29] = 1'b0;
    assign proc_7_data_PIPO_blk[29] = 1'b0;
    assign proc_7_start_FIFO_blk[29] = 1'b0;
    assign proc_7_TLF_FIFO_blk[29] = 1'b0;
    assign proc_7_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_7_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_7[29] = dl_detect_out ? proc_dep_vld_vec_7_reg[29] : (proc_7_data_FIFO_blk[29] | proc_7_data_PIPO_blk[29] | proc_7_start_FIFO_blk[29] | proc_7_TLF_FIFO_blk[29] | proc_7_input_sync_blk[29] | proc_7_output_sync_blk[29]);
    assign proc_7_data_FIFO_blk[30] = 1'b0;
    assign proc_7_data_PIPO_blk[30] = 1'b0;
    assign proc_7_start_FIFO_blk[30] = 1'b0;
    assign proc_7_TLF_FIFO_blk[30] = 1'b0;
    assign proc_7_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_7_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_7[30] = dl_detect_out ? proc_dep_vld_vec_7_reg[30] : (proc_7_data_FIFO_blk[30] | proc_7_data_PIPO_blk[30] | proc_7_start_FIFO_blk[30] | proc_7_TLF_FIFO_blk[30] | proc_7_input_sync_blk[30] | proc_7_output_sync_blk[30]);
    assign proc_7_data_FIFO_blk[31] = 1'b0;
    assign proc_7_data_PIPO_blk[31] = 1'b0;
    assign proc_7_start_FIFO_blk[31] = 1'b0;
    assign proc_7_TLF_FIFO_blk[31] = 1'b0;
    assign proc_7_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_7_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_7[31] = dl_detect_out ? proc_dep_vld_vec_7_reg[31] : (proc_7_data_FIFO_blk[31] | proc_7_data_PIPO_blk[31] | proc_7_start_FIFO_blk[31] | proc_7_TLF_FIFO_blk[31] | proc_7_input_sync_blk[31] | proc_7_output_sync_blk[31]);
    assign proc_7_data_FIFO_blk[32] = 1'b0;
    assign proc_7_data_PIPO_blk[32] = 1'b0;
    assign proc_7_start_FIFO_blk[32] = 1'b0;
    assign proc_7_TLF_FIFO_blk[32] = 1'b0;
    assign proc_7_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_2_U0_ap_ready & ProcessingElement_2_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_7_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_7[32] = dl_detect_out ? proc_dep_vld_vec_7_reg[32] : (proc_7_data_FIFO_blk[32] | proc_7_data_PIPO_blk[32] | proc_7_start_FIFO_blk[32] | proc_7_TLF_FIFO_blk[32] | proc_7_input_sync_blk[32] | proc_7_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_7_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_7_reg <= proc_dep_vld_vec_7;
        end
    end
    assign in_chan_dep_vld_vec_7[0] = dep_chan_vld_0_7;
    assign in_chan_dep_data_vec_7[39 : 0] = dep_chan_data_0_7;
    assign token_in_vec_7[0] = token_0_7;
    assign in_chan_dep_vld_vec_7[1] = dep_chan_vld_1_7;
    assign in_chan_dep_data_vec_7[79 : 40] = dep_chan_data_1_7;
    assign token_in_vec_7[1] = token_1_7;
    assign in_chan_dep_vld_vec_7[2] = dep_chan_vld_3_7;
    assign in_chan_dep_data_vec_7[119 : 80] = dep_chan_data_3_7;
    assign token_in_vec_7[2] = token_3_7;
    assign in_chan_dep_vld_vec_7[3] = dep_chan_vld_6_7;
    assign in_chan_dep_data_vec_7[159 : 120] = dep_chan_data_6_7;
    assign token_in_vec_7[3] = token_6_7;
    assign in_chan_dep_vld_vec_7[4] = dep_chan_vld_8_7;
    assign in_chan_dep_data_vec_7[199 : 160] = dep_chan_data_8_7;
    assign token_in_vec_7[4] = token_8_7;
    assign in_chan_dep_vld_vec_7[5] = dep_chan_vld_9_7;
    assign in_chan_dep_data_vec_7[239 : 200] = dep_chan_data_9_7;
    assign token_in_vec_7[5] = token_9_7;
    assign in_chan_dep_vld_vec_7[6] = dep_chan_vld_10_7;
    assign in_chan_dep_data_vec_7[279 : 240] = dep_chan_data_10_7;
    assign token_in_vec_7[6] = token_10_7;
    assign in_chan_dep_vld_vec_7[7] = dep_chan_vld_11_7;
    assign in_chan_dep_data_vec_7[319 : 280] = dep_chan_data_11_7;
    assign token_in_vec_7[7] = token_11_7;
    assign in_chan_dep_vld_vec_7[8] = dep_chan_vld_12_7;
    assign in_chan_dep_data_vec_7[359 : 320] = dep_chan_data_12_7;
    assign token_in_vec_7[8] = token_12_7;
    assign in_chan_dep_vld_vec_7[9] = dep_chan_vld_13_7;
    assign in_chan_dep_data_vec_7[399 : 360] = dep_chan_data_13_7;
    assign token_in_vec_7[9] = token_13_7;
    assign in_chan_dep_vld_vec_7[10] = dep_chan_vld_14_7;
    assign in_chan_dep_data_vec_7[439 : 400] = dep_chan_data_14_7;
    assign token_in_vec_7[10] = token_14_7;
    assign in_chan_dep_vld_vec_7[11] = dep_chan_vld_15_7;
    assign in_chan_dep_data_vec_7[479 : 440] = dep_chan_data_15_7;
    assign token_in_vec_7[11] = token_15_7;
    assign in_chan_dep_vld_vec_7[12] = dep_chan_vld_16_7;
    assign in_chan_dep_data_vec_7[519 : 480] = dep_chan_data_16_7;
    assign token_in_vec_7[12] = token_16_7;
    assign in_chan_dep_vld_vec_7[13] = dep_chan_vld_17_7;
    assign in_chan_dep_data_vec_7[559 : 520] = dep_chan_data_17_7;
    assign token_in_vec_7[13] = token_17_7;
    assign in_chan_dep_vld_vec_7[14] = dep_chan_vld_18_7;
    assign in_chan_dep_data_vec_7[599 : 560] = dep_chan_data_18_7;
    assign token_in_vec_7[14] = token_18_7;
    assign in_chan_dep_vld_vec_7[15] = dep_chan_vld_19_7;
    assign in_chan_dep_data_vec_7[639 : 600] = dep_chan_data_19_7;
    assign token_in_vec_7[15] = token_19_7;
    assign in_chan_dep_vld_vec_7[16] = dep_chan_vld_20_7;
    assign in_chan_dep_data_vec_7[679 : 640] = dep_chan_data_20_7;
    assign token_in_vec_7[16] = token_20_7;
    assign in_chan_dep_vld_vec_7[17] = dep_chan_vld_21_7;
    assign in_chan_dep_data_vec_7[719 : 680] = dep_chan_data_21_7;
    assign token_in_vec_7[17] = token_21_7;
    assign in_chan_dep_vld_vec_7[18] = dep_chan_vld_22_7;
    assign in_chan_dep_data_vec_7[759 : 720] = dep_chan_data_22_7;
    assign token_in_vec_7[18] = token_22_7;
    assign in_chan_dep_vld_vec_7[19] = dep_chan_vld_23_7;
    assign in_chan_dep_data_vec_7[799 : 760] = dep_chan_data_23_7;
    assign token_in_vec_7[19] = token_23_7;
    assign in_chan_dep_vld_vec_7[20] = dep_chan_vld_24_7;
    assign in_chan_dep_data_vec_7[839 : 800] = dep_chan_data_24_7;
    assign token_in_vec_7[20] = token_24_7;
    assign in_chan_dep_vld_vec_7[21] = dep_chan_vld_25_7;
    assign in_chan_dep_data_vec_7[879 : 840] = dep_chan_data_25_7;
    assign token_in_vec_7[21] = token_25_7;
    assign in_chan_dep_vld_vec_7[22] = dep_chan_vld_26_7;
    assign in_chan_dep_data_vec_7[919 : 880] = dep_chan_data_26_7;
    assign token_in_vec_7[22] = token_26_7;
    assign in_chan_dep_vld_vec_7[23] = dep_chan_vld_27_7;
    assign in_chan_dep_data_vec_7[959 : 920] = dep_chan_data_27_7;
    assign token_in_vec_7[23] = token_27_7;
    assign in_chan_dep_vld_vec_7[24] = dep_chan_vld_28_7;
    assign in_chan_dep_data_vec_7[999 : 960] = dep_chan_data_28_7;
    assign token_in_vec_7[24] = token_28_7;
    assign in_chan_dep_vld_vec_7[25] = dep_chan_vld_29_7;
    assign in_chan_dep_data_vec_7[1039 : 1000] = dep_chan_data_29_7;
    assign token_in_vec_7[25] = token_29_7;
    assign in_chan_dep_vld_vec_7[26] = dep_chan_vld_30_7;
    assign in_chan_dep_data_vec_7[1079 : 1040] = dep_chan_data_30_7;
    assign token_in_vec_7[26] = token_30_7;
    assign in_chan_dep_vld_vec_7[27] = dep_chan_vld_31_7;
    assign in_chan_dep_data_vec_7[1119 : 1080] = dep_chan_data_31_7;
    assign token_in_vec_7[27] = token_31_7;
    assign in_chan_dep_vld_vec_7[28] = dep_chan_vld_32_7;
    assign in_chan_dep_data_vec_7[1159 : 1120] = dep_chan_data_32_7;
    assign token_in_vec_7[28] = token_32_7;
    assign in_chan_dep_vld_vec_7[29] = dep_chan_vld_33_7;
    assign in_chan_dep_data_vec_7[1199 : 1160] = dep_chan_data_33_7;
    assign token_in_vec_7[29] = token_33_7;
    assign in_chan_dep_vld_vec_7[30] = dep_chan_vld_34_7;
    assign in_chan_dep_data_vec_7[1239 : 1200] = dep_chan_data_34_7;
    assign token_in_vec_7[30] = token_34_7;
    assign in_chan_dep_vld_vec_7[31] = dep_chan_vld_35_7;
    assign in_chan_dep_data_vec_7[1279 : 1240] = dep_chan_data_35_7;
    assign token_in_vec_7[31] = token_35_7;
    assign in_chan_dep_vld_vec_7[32] = dep_chan_vld_36_7;
    assign in_chan_dep_data_vec_7[1319 : 1280] = dep_chan_data_36_7;
    assign token_in_vec_7[32] = token_36_7;
    assign dep_chan_vld_7_6 = out_chan_dep_vld_vec_7[0];
    assign dep_chan_data_7_6 = out_chan_dep_data_7;
    assign token_7_6 = token_out_vec_7[0];
    assign dep_chan_vld_7_8 = out_chan_dep_vld_vec_7[1];
    assign dep_chan_data_7_8 = out_chan_dep_data_7;
    assign token_7_8 = token_out_vec_7[1];
    assign dep_chan_vld_7_0 = out_chan_dep_vld_vec_7[2];
    assign dep_chan_data_7_0 = out_chan_dep_data_7;
    assign token_7_0 = token_out_vec_7[2];
    assign dep_chan_vld_7_1 = out_chan_dep_vld_vec_7[3];
    assign dep_chan_data_7_1 = out_chan_dep_data_7;
    assign token_7_1 = token_out_vec_7[3];
    assign dep_chan_vld_7_3 = out_chan_dep_vld_vec_7[4];
    assign dep_chan_data_7_3 = out_chan_dep_data_7;
    assign token_7_3 = token_out_vec_7[4];
    assign dep_chan_vld_7_9 = out_chan_dep_vld_vec_7[5];
    assign dep_chan_data_7_9 = out_chan_dep_data_7;
    assign token_7_9 = token_out_vec_7[5];
    assign dep_chan_vld_7_10 = out_chan_dep_vld_vec_7[6];
    assign dep_chan_data_7_10 = out_chan_dep_data_7;
    assign token_7_10 = token_out_vec_7[6];
    assign dep_chan_vld_7_11 = out_chan_dep_vld_vec_7[7];
    assign dep_chan_data_7_11 = out_chan_dep_data_7;
    assign token_7_11 = token_out_vec_7[7];
    assign dep_chan_vld_7_12 = out_chan_dep_vld_vec_7[8];
    assign dep_chan_data_7_12 = out_chan_dep_data_7;
    assign token_7_12 = token_out_vec_7[8];
    assign dep_chan_vld_7_13 = out_chan_dep_vld_vec_7[9];
    assign dep_chan_data_7_13 = out_chan_dep_data_7;
    assign token_7_13 = token_out_vec_7[9];
    assign dep_chan_vld_7_14 = out_chan_dep_vld_vec_7[10];
    assign dep_chan_data_7_14 = out_chan_dep_data_7;
    assign token_7_14 = token_out_vec_7[10];
    assign dep_chan_vld_7_15 = out_chan_dep_vld_vec_7[11];
    assign dep_chan_data_7_15 = out_chan_dep_data_7;
    assign token_7_15 = token_out_vec_7[11];
    assign dep_chan_vld_7_16 = out_chan_dep_vld_vec_7[12];
    assign dep_chan_data_7_16 = out_chan_dep_data_7;
    assign token_7_16 = token_out_vec_7[12];
    assign dep_chan_vld_7_17 = out_chan_dep_vld_vec_7[13];
    assign dep_chan_data_7_17 = out_chan_dep_data_7;
    assign token_7_17 = token_out_vec_7[13];
    assign dep_chan_vld_7_18 = out_chan_dep_vld_vec_7[14];
    assign dep_chan_data_7_18 = out_chan_dep_data_7;
    assign token_7_18 = token_out_vec_7[14];
    assign dep_chan_vld_7_19 = out_chan_dep_vld_vec_7[15];
    assign dep_chan_data_7_19 = out_chan_dep_data_7;
    assign token_7_19 = token_out_vec_7[15];
    assign dep_chan_vld_7_20 = out_chan_dep_vld_vec_7[16];
    assign dep_chan_data_7_20 = out_chan_dep_data_7;
    assign token_7_20 = token_out_vec_7[16];
    assign dep_chan_vld_7_21 = out_chan_dep_vld_vec_7[17];
    assign dep_chan_data_7_21 = out_chan_dep_data_7;
    assign token_7_21 = token_out_vec_7[17];
    assign dep_chan_vld_7_22 = out_chan_dep_vld_vec_7[18];
    assign dep_chan_data_7_22 = out_chan_dep_data_7;
    assign token_7_22 = token_out_vec_7[18];
    assign dep_chan_vld_7_23 = out_chan_dep_vld_vec_7[19];
    assign dep_chan_data_7_23 = out_chan_dep_data_7;
    assign token_7_23 = token_out_vec_7[19];
    assign dep_chan_vld_7_24 = out_chan_dep_vld_vec_7[20];
    assign dep_chan_data_7_24 = out_chan_dep_data_7;
    assign token_7_24 = token_out_vec_7[20];
    assign dep_chan_vld_7_25 = out_chan_dep_vld_vec_7[21];
    assign dep_chan_data_7_25 = out_chan_dep_data_7;
    assign token_7_25 = token_out_vec_7[21];
    assign dep_chan_vld_7_26 = out_chan_dep_vld_vec_7[22];
    assign dep_chan_data_7_26 = out_chan_dep_data_7;
    assign token_7_26 = token_out_vec_7[22];
    assign dep_chan_vld_7_27 = out_chan_dep_vld_vec_7[23];
    assign dep_chan_data_7_27 = out_chan_dep_data_7;
    assign token_7_27 = token_out_vec_7[23];
    assign dep_chan_vld_7_28 = out_chan_dep_vld_vec_7[24];
    assign dep_chan_data_7_28 = out_chan_dep_data_7;
    assign token_7_28 = token_out_vec_7[24];
    assign dep_chan_vld_7_29 = out_chan_dep_vld_vec_7[25];
    assign dep_chan_data_7_29 = out_chan_dep_data_7;
    assign token_7_29 = token_out_vec_7[25];
    assign dep_chan_vld_7_30 = out_chan_dep_vld_vec_7[26];
    assign dep_chan_data_7_30 = out_chan_dep_data_7;
    assign token_7_30 = token_out_vec_7[26];
    assign dep_chan_vld_7_31 = out_chan_dep_vld_vec_7[27];
    assign dep_chan_data_7_31 = out_chan_dep_data_7;
    assign token_7_31 = token_out_vec_7[27];
    assign dep_chan_vld_7_32 = out_chan_dep_vld_vec_7[28];
    assign dep_chan_data_7_32 = out_chan_dep_data_7;
    assign token_7_32 = token_out_vec_7[28];
    assign dep_chan_vld_7_33 = out_chan_dep_vld_vec_7[29];
    assign dep_chan_data_7_33 = out_chan_dep_data_7;
    assign token_7_33 = token_out_vec_7[29];
    assign dep_chan_vld_7_34 = out_chan_dep_vld_vec_7[30];
    assign dep_chan_data_7_34 = out_chan_dep_data_7;
    assign token_7_34 = token_out_vec_7[30];
    assign dep_chan_vld_7_35 = out_chan_dep_vld_vec_7[31];
    assign dep_chan_data_7_35 = out_chan_dep_data_7;
    assign token_7_35 = token_out_vec_7[31];
    assign dep_chan_vld_7_36 = out_chan_dep_vld_vec_7[32];
    assign dep_chan_data_7_36 = out_chan_dep_data_7;
    assign token_7_36 = token_out_vec_7[32];

    // Process: ProcessingElement_3_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 8, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_8 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_8),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_8),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_8),
        .token_in_vec(token_in_vec_8),
        .dl_detect_in(dl_detect_out),
        .origin(origin[8]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_8),
        .out_chan_dep_data(out_chan_dep_data_8),
        .token_out_vec(token_out_vec_8),
        .dl_detect_out(dl_in_vec[8]));

    assign proc_8_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_2_blk_n) | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_2_blk_n) | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_WriteC_Flattened_fu_179.cPipes_2_blk_n);
    assign proc_8_data_PIPO_blk[0] = 1'b0;
    assign proc_8_start_FIFO_blk[0] = 1'b0;
    assign proc_8_TLF_FIFO_blk[0] = 1'b0;
    assign proc_8_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_8_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_8[0] = dl_detect_out ? proc_dep_vld_vec_8_reg[0] : (proc_8_data_FIFO_blk[0] | proc_8_data_PIPO_blk[0] | proc_8_start_FIFO_blk[0] | proc_8_TLF_FIFO_blk[0] | proc_8_input_sync_blk[0] | proc_8_output_sync_blk[0]);
    assign proc_8_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_3_blk_n) | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_3_blk_n) | (~ProcessingElement_3_U0.grp_ProcessingElement_3_Pipeline_WriteC_Flattened_fu_179.cPipes_3_blk_n);
    assign proc_8_data_PIPO_blk[1] = 1'b0;
    assign proc_8_start_FIFO_blk[1] = 1'b0;
    assign proc_8_TLF_FIFO_blk[1] = 1'b0;
    assign proc_8_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_8_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_8[1] = dl_detect_out ? proc_dep_vld_vec_8_reg[1] : (proc_8_data_FIFO_blk[1] | proc_8_data_PIPO_blk[1] | proc_8_start_FIFO_blk[1] | proc_8_TLF_FIFO_blk[1] | proc_8_input_sync_blk[1] | proc_8_output_sync_blk[1]);
    assign proc_8_data_FIFO_blk[2] = 1'b0;
    assign proc_8_data_PIPO_blk[2] = 1'b0;
    assign proc_8_start_FIFO_blk[2] = 1'b0;
    assign proc_8_TLF_FIFO_blk[2] = 1'b0;
    assign proc_8_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_8_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_8[2] = dl_detect_out ? proc_dep_vld_vec_8_reg[2] : (proc_8_data_FIFO_blk[2] | proc_8_data_PIPO_blk[2] | proc_8_start_FIFO_blk[2] | proc_8_TLF_FIFO_blk[2] | proc_8_input_sync_blk[2] | proc_8_output_sync_blk[2]);
    assign proc_8_data_FIFO_blk[3] = 1'b0;
    assign proc_8_data_PIPO_blk[3] = 1'b0;
    assign proc_8_start_FIFO_blk[3] = 1'b0;
    assign proc_8_TLF_FIFO_blk[3] = 1'b0;
    assign proc_8_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_8_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_8[3] = dl_detect_out ? proc_dep_vld_vec_8_reg[3] : (proc_8_data_FIFO_blk[3] | proc_8_data_PIPO_blk[3] | proc_8_start_FIFO_blk[3] | proc_8_TLF_FIFO_blk[3] | proc_8_input_sync_blk[3] | proc_8_output_sync_blk[3]);
    assign proc_8_data_FIFO_blk[4] = 1'b0;
    assign proc_8_data_PIPO_blk[4] = 1'b0;
    assign proc_8_start_FIFO_blk[4] = 1'b0;
    assign proc_8_TLF_FIFO_blk[4] = 1'b0;
    assign proc_8_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_8_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_8[4] = dl_detect_out ? proc_dep_vld_vec_8_reg[4] : (proc_8_data_FIFO_blk[4] | proc_8_data_PIPO_blk[4] | proc_8_start_FIFO_blk[4] | proc_8_TLF_FIFO_blk[4] | proc_8_input_sync_blk[4] | proc_8_output_sync_blk[4]);
    assign proc_8_data_FIFO_blk[5] = 1'b0;
    assign proc_8_data_PIPO_blk[5] = 1'b0;
    assign proc_8_start_FIFO_blk[5] = 1'b0;
    assign proc_8_TLF_FIFO_blk[5] = 1'b0;
    assign proc_8_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_8_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_8[5] = dl_detect_out ? proc_dep_vld_vec_8_reg[5] : (proc_8_data_FIFO_blk[5] | proc_8_data_PIPO_blk[5] | proc_8_start_FIFO_blk[5] | proc_8_TLF_FIFO_blk[5] | proc_8_input_sync_blk[5] | proc_8_output_sync_blk[5]);
    assign proc_8_data_FIFO_blk[6] = 1'b0;
    assign proc_8_data_PIPO_blk[6] = 1'b0;
    assign proc_8_start_FIFO_blk[6] = 1'b0;
    assign proc_8_TLF_FIFO_blk[6] = 1'b0;
    assign proc_8_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_8_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_8[6] = dl_detect_out ? proc_dep_vld_vec_8_reg[6] : (proc_8_data_FIFO_blk[6] | proc_8_data_PIPO_blk[6] | proc_8_start_FIFO_blk[6] | proc_8_TLF_FIFO_blk[6] | proc_8_input_sync_blk[6] | proc_8_output_sync_blk[6]);
    assign proc_8_data_FIFO_blk[7] = 1'b0;
    assign proc_8_data_PIPO_blk[7] = 1'b0;
    assign proc_8_start_FIFO_blk[7] = 1'b0;
    assign proc_8_TLF_FIFO_blk[7] = 1'b0;
    assign proc_8_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_8_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_8[7] = dl_detect_out ? proc_dep_vld_vec_8_reg[7] : (proc_8_data_FIFO_blk[7] | proc_8_data_PIPO_blk[7] | proc_8_start_FIFO_blk[7] | proc_8_TLF_FIFO_blk[7] | proc_8_input_sync_blk[7] | proc_8_output_sync_blk[7]);
    assign proc_8_data_FIFO_blk[8] = 1'b0;
    assign proc_8_data_PIPO_blk[8] = 1'b0;
    assign proc_8_start_FIFO_blk[8] = 1'b0;
    assign proc_8_TLF_FIFO_blk[8] = 1'b0;
    assign proc_8_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_8_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_8[8] = dl_detect_out ? proc_dep_vld_vec_8_reg[8] : (proc_8_data_FIFO_blk[8] | proc_8_data_PIPO_blk[8] | proc_8_start_FIFO_blk[8] | proc_8_TLF_FIFO_blk[8] | proc_8_input_sync_blk[8] | proc_8_output_sync_blk[8]);
    assign proc_8_data_FIFO_blk[9] = 1'b0;
    assign proc_8_data_PIPO_blk[9] = 1'b0;
    assign proc_8_start_FIFO_blk[9] = 1'b0;
    assign proc_8_TLF_FIFO_blk[9] = 1'b0;
    assign proc_8_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_8_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_8[9] = dl_detect_out ? proc_dep_vld_vec_8_reg[9] : (proc_8_data_FIFO_blk[9] | proc_8_data_PIPO_blk[9] | proc_8_start_FIFO_blk[9] | proc_8_TLF_FIFO_blk[9] | proc_8_input_sync_blk[9] | proc_8_output_sync_blk[9]);
    assign proc_8_data_FIFO_blk[10] = 1'b0;
    assign proc_8_data_PIPO_blk[10] = 1'b0;
    assign proc_8_start_FIFO_blk[10] = 1'b0;
    assign proc_8_TLF_FIFO_blk[10] = 1'b0;
    assign proc_8_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_8_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_8[10] = dl_detect_out ? proc_dep_vld_vec_8_reg[10] : (proc_8_data_FIFO_blk[10] | proc_8_data_PIPO_blk[10] | proc_8_start_FIFO_blk[10] | proc_8_TLF_FIFO_blk[10] | proc_8_input_sync_blk[10] | proc_8_output_sync_blk[10]);
    assign proc_8_data_FIFO_blk[11] = 1'b0;
    assign proc_8_data_PIPO_blk[11] = 1'b0;
    assign proc_8_start_FIFO_blk[11] = 1'b0;
    assign proc_8_TLF_FIFO_blk[11] = 1'b0;
    assign proc_8_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_8_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_8[11] = dl_detect_out ? proc_dep_vld_vec_8_reg[11] : (proc_8_data_FIFO_blk[11] | proc_8_data_PIPO_blk[11] | proc_8_start_FIFO_blk[11] | proc_8_TLF_FIFO_blk[11] | proc_8_input_sync_blk[11] | proc_8_output_sync_blk[11]);
    assign proc_8_data_FIFO_blk[12] = 1'b0;
    assign proc_8_data_PIPO_blk[12] = 1'b0;
    assign proc_8_start_FIFO_blk[12] = 1'b0;
    assign proc_8_TLF_FIFO_blk[12] = 1'b0;
    assign proc_8_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_8_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_8[12] = dl_detect_out ? proc_dep_vld_vec_8_reg[12] : (proc_8_data_FIFO_blk[12] | proc_8_data_PIPO_blk[12] | proc_8_start_FIFO_blk[12] | proc_8_TLF_FIFO_blk[12] | proc_8_input_sync_blk[12] | proc_8_output_sync_blk[12]);
    assign proc_8_data_FIFO_blk[13] = 1'b0;
    assign proc_8_data_PIPO_blk[13] = 1'b0;
    assign proc_8_start_FIFO_blk[13] = 1'b0;
    assign proc_8_TLF_FIFO_blk[13] = 1'b0;
    assign proc_8_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_8_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_8[13] = dl_detect_out ? proc_dep_vld_vec_8_reg[13] : (proc_8_data_FIFO_blk[13] | proc_8_data_PIPO_blk[13] | proc_8_start_FIFO_blk[13] | proc_8_TLF_FIFO_blk[13] | proc_8_input_sync_blk[13] | proc_8_output_sync_blk[13]);
    assign proc_8_data_FIFO_blk[14] = 1'b0;
    assign proc_8_data_PIPO_blk[14] = 1'b0;
    assign proc_8_start_FIFO_blk[14] = 1'b0;
    assign proc_8_TLF_FIFO_blk[14] = 1'b0;
    assign proc_8_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_8_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_8[14] = dl_detect_out ? proc_dep_vld_vec_8_reg[14] : (proc_8_data_FIFO_blk[14] | proc_8_data_PIPO_blk[14] | proc_8_start_FIFO_blk[14] | proc_8_TLF_FIFO_blk[14] | proc_8_input_sync_blk[14] | proc_8_output_sync_blk[14]);
    assign proc_8_data_FIFO_blk[15] = 1'b0;
    assign proc_8_data_PIPO_blk[15] = 1'b0;
    assign proc_8_start_FIFO_blk[15] = 1'b0;
    assign proc_8_TLF_FIFO_blk[15] = 1'b0;
    assign proc_8_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_8_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_8[15] = dl_detect_out ? proc_dep_vld_vec_8_reg[15] : (proc_8_data_FIFO_blk[15] | proc_8_data_PIPO_blk[15] | proc_8_start_FIFO_blk[15] | proc_8_TLF_FIFO_blk[15] | proc_8_input_sync_blk[15] | proc_8_output_sync_blk[15]);
    assign proc_8_data_FIFO_blk[16] = 1'b0;
    assign proc_8_data_PIPO_blk[16] = 1'b0;
    assign proc_8_start_FIFO_blk[16] = 1'b0;
    assign proc_8_TLF_FIFO_blk[16] = 1'b0;
    assign proc_8_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_8_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_8[16] = dl_detect_out ? proc_dep_vld_vec_8_reg[16] : (proc_8_data_FIFO_blk[16] | proc_8_data_PIPO_blk[16] | proc_8_start_FIFO_blk[16] | proc_8_TLF_FIFO_blk[16] | proc_8_input_sync_blk[16] | proc_8_output_sync_blk[16]);
    assign proc_8_data_FIFO_blk[17] = 1'b0;
    assign proc_8_data_PIPO_blk[17] = 1'b0;
    assign proc_8_start_FIFO_blk[17] = 1'b0;
    assign proc_8_TLF_FIFO_blk[17] = 1'b0;
    assign proc_8_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_8_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_8[17] = dl_detect_out ? proc_dep_vld_vec_8_reg[17] : (proc_8_data_FIFO_blk[17] | proc_8_data_PIPO_blk[17] | proc_8_start_FIFO_blk[17] | proc_8_TLF_FIFO_blk[17] | proc_8_input_sync_blk[17] | proc_8_output_sync_blk[17]);
    assign proc_8_data_FIFO_blk[18] = 1'b0;
    assign proc_8_data_PIPO_blk[18] = 1'b0;
    assign proc_8_start_FIFO_blk[18] = 1'b0;
    assign proc_8_TLF_FIFO_blk[18] = 1'b0;
    assign proc_8_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_8_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_8[18] = dl_detect_out ? proc_dep_vld_vec_8_reg[18] : (proc_8_data_FIFO_blk[18] | proc_8_data_PIPO_blk[18] | proc_8_start_FIFO_blk[18] | proc_8_TLF_FIFO_blk[18] | proc_8_input_sync_blk[18] | proc_8_output_sync_blk[18]);
    assign proc_8_data_FIFO_blk[19] = 1'b0;
    assign proc_8_data_PIPO_blk[19] = 1'b0;
    assign proc_8_start_FIFO_blk[19] = 1'b0;
    assign proc_8_TLF_FIFO_blk[19] = 1'b0;
    assign proc_8_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_8_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_8[19] = dl_detect_out ? proc_dep_vld_vec_8_reg[19] : (proc_8_data_FIFO_blk[19] | proc_8_data_PIPO_blk[19] | proc_8_start_FIFO_blk[19] | proc_8_TLF_FIFO_blk[19] | proc_8_input_sync_blk[19] | proc_8_output_sync_blk[19]);
    assign proc_8_data_FIFO_blk[20] = 1'b0;
    assign proc_8_data_PIPO_blk[20] = 1'b0;
    assign proc_8_start_FIFO_blk[20] = 1'b0;
    assign proc_8_TLF_FIFO_blk[20] = 1'b0;
    assign proc_8_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_8_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_8[20] = dl_detect_out ? proc_dep_vld_vec_8_reg[20] : (proc_8_data_FIFO_blk[20] | proc_8_data_PIPO_blk[20] | proc_8_start_FIFO_blk[20] | proc_8_TLF_FIFO_blk[20] | proc_8_input_sync_blk[20] | proc_8_output_sync_blk[20]);
    assign proc_8_data_FIFO_blk[21] = 1'b0;
    assign proc_8_data_PIPO_blk[21] = 1'b0;
    assign proc_8_start_FIFO_blk[21] = 1'b0;
    assign proc_8_TLF_FIFO_blk[21] = 1'b0;
    assign proc_8_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_8_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_8[21] = dl_detect_out ? proc_dep_vld_vec_8_reg[21] : (proc_8_data_FIFO_blk[21] | proc_8_data_PIPO_blk[21] | proc_8_start_FIFO_blk[21] | proc_8_TLF_FIFO_blk[21] | proc_8_input_sync_blk[21] | proc_8_output_sync_blk[21]);
    assign proc_8_data_FIFO_blk[22] = 1'b0;
    assign proc_8_data_PIPO_blk[22] = 1'b0;
    assign proc_8_start_FIFO_blk[22] = 1'b0;
    assign proc_8_TLF_FIFO_blk[22] = 1'b0;
    assign proc_8_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_8_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_8[22] = dl_detect_out ? proc_dep_vld_vec_8_reg[22] : (proc_8_data_FIFO_blk[22] | proc_8_data_PIPO_blk[22] | proc_8_start_FIFO_blk[22] | proc_8_TLF_FIFO_blk[22] | proc_8_input_sync_blk[22] | proc_8_output_sync_blk[22]);
    assign proc_8_data_FIFO_blk[23] = 1'b0;
    assign proc_8_data_PIPO_blk[23] = 1'b0;
    assign proc_8_start_FIFO_blk[23] = 1'b0;
    assign proc_8_TLF_FIFO_blk[23] = 1'b0;
    assign proc_8_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_8_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_8[23] = dl_detect_out ? proc_dep_vld_vec_8_reg[23] : (proc_8_data_FIFO_blk[23] | proc_8_data_PIPO_blk[23] | proc_8_start_FIFO_blk[23] | proc_8_TLF_FIFO_blk[23] | proc_8_input_sync_blk[23] | proc_8_output_sync_blk[23]);
    assign proc_8_data_FIFO_blk[24] = 1'b0;
    assign proc_8_data_PIPO_blk[24] = 1'b0;
    assign proc_8_start_FIFO_blk[24] = 1'b0;
    assign proc_8_TLF_FIFO_blk[24] = 1'b0;
    assign proc_8_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_8_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_8[24] = dl_detect_out ? proc_dep_vld_vec_8_reg[24] : (proc_8_data_FIFO_blk[24] | proc_8_data_PIPO_blk[24] | proc_8_start_FIFO_blk[24] | proc_8_TLF_FIFO_blk[24] | proc_8_input_sync_blk[24] | proc_8_output_sync_blk[24]);
    assign proc_8_data_FIFO_blk[25] = 1'b0;
    assign proc_8_data_PIPO_blk[25] = 1'b0;
    assign proc_8_start_FIFO_blk[25] = 1'b0;
    assign proc_8_TLF_FIFO_blk[25] = 1'b0;
    assign proc_8_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_8_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_8[25] = dl_detect_out ? proc_dep_vld_vec_8_reg[25] : (proc_8_data_FIFO_blk[25] | proc_8_data_PIPO_blk[25] | proc_8_start_FIFO_blk[25] | proc_8_TLF_FIFO_blk[25] | proc_8_input_sync_blk[25] | proc_8_output_sync_blk[25]);
    assign proc_8_data_FIFO_blk[26] = 1'b0;
    assign proc_8_data_PIPO_blk[26] = 1'b0;
    assign proc_8_start_FIFO_blk[26] = 1'b0;
    assign proc_8_TLF_FIFO_blk[26] = 1'b0;
    assign proc_8_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_8_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_8[26] = dl_detect_out ? proc_dep_vld_vec_8_reg[26] : (proc_8_data_FIFO_blk[26] | proc_8_data_PIPO_blk[26] | proc_8_start_FIFO_blk[26] | proc_8_TLF_FIFO_blk[26] | proc_8_input_sync_blk[26] | proc_8_output_sync_blk[26]);
    assign proc_8_data_FIFO_blk[27] = 1'b0;
    assign proc_8_data_PIPO_blk[27] = 1'b0;
    assign proc_8_start_FIFO_blk[27] = 1'b0;
    assign proc_8_TLF_FIFO_blk[27] = 1'b0;
    assign proc_8_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_8_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_8[27] = dl_detect_out ? proc_dep_vld_vec_8_reg[27] : (proc_8_data_FIFO_blk[27] | proc_8_data_PIPO_blk[27] | proc_8_start_FIFO_blk[27] | proc_8_TLF_FIFO_blk[27] | proc_8_input_sync_blk[27] | proc_8_output_sync_blk[27]);
    assign proc_8_data_FIFO_blk[28] = 1'b0;
    assign proc_8_data_PIPO_blk[28] = 1'b0;
    assign proc_8_start_FIFO_blk[28] = 1'b0;
    assign proc_8_TLF_FIFO_blk[28] = 1'b0;
    assign proc_8_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_8_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_8[28] = dl_detect_out ? proc_dep_vld_vec_8_reg[28] : (proc_8_data_FIFO_blk[28] | proc_8_data_PIPO_blk[28] | proc_8_start_FIFO_blk[28] | proc_8_TLF_FIFO_blk[28] | proc_8_input_sync_blk[28] | proc_8_output_sync_blk[28]);
    assign proc_8_data_FIFO_blk[29] = 1'b0;
    assign proc_8_data_PIPO_blk[29] = 1'b0;
    assign proc_8_start_FIFO_blk[29] = 1'b0;
    assign proc_8_TLF_FIFO_blk[29] = 1'b0;
    assign proc_8_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_8_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_8[29] = dl_detect_out ? proc_dep_vld_vec_8_reg[29] : (proc_8_data_FIFO_blk[29] | proc_8_data_PIPO_blk[29] | proc_8_start_FIFO_blk[29] | proc_8_TLF_FIFO_blk[29] | proc_8_input_sync_blk[29] | proc_8_output_sync_blk[29]);
    assign proc_8_data_FIFO_blk[30] = 1'b0;
    assign proc_8_data_PIPO_blk[30] = 1'b0;
    assign proc_8_start_FIFO_blk[30] = 1'b0;
    assign proc_8_TLF_FIFO_blk[30] = 1'b0;
    assign proc_8_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_8_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_8[30] = dl_detect_out ? proc_dep_vld_vec_8_reg[30] : (proc_8_data_FIFO_blk[30] | proc_8_data_PIPO_blk[30] | proc_8_start_FIFO_blk[30] | proc_8_TLF_FIFO_blk[30] | proc_8_input_sync_blk[30] | proc_8_output_sync_blk[30]);
    assign proc_8_data_FIFO_blk[31] = 1'b0;
    assign proc_8_data_PIPO_blk[31] = 1'b0;
    assign proc_8_start_FIFO_blk[31] = 1'b0;
    assign proc_8_TLF_FIFO_blk[31] = 1'b0;
    assign proc_8_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_8_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_8[31] = dl_detect_out ? proc_dep_vld_vec_8_reg[31] : (proc_8_data_FIFO_blk[31] | proc_8_data_PIPO_blk[31] | proc_8_start_FIFO_blk[31] | proc_8_TLF_FIFO_blk[31] | proc_8_input_sync_blk[31] | proc_8_output_sync_blk[31]);
    assign proc_8_data_FIFO_blk[32] = 1'b0;
    assign proc_8_data_PIPO_blk[32] = 1'b0;
    assign proc_8_start_FIFO_blk[32] = 1'b0;
    assign proc_8_TLF_FIFO_blk[32] = 1'b0;
    assign proc_8_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_3_U0_ap_ready & ProcessingElement_3_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_8_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_8[32] = dl_detect_out ? proc_dep_vld_vec_8_reg[32] : (proc_8_data_FIFO_blk[32] | proc_8_data_PIPO_blk[32] | proc_8_start_FIFO_blk[32] | proc_8_TLF_FIFO_blk[32] | proc_8_input_sync_blk[32] | proc_8_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_8_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_8_reg <= proc_dep_vld_vec_8;
        end
    end
    assign in_chan_dep_vld_vec_8[0] = dep_chan_vld_0_8;
    assign in_chan_dep_data_vec_8[39 : 0] = dep_chan_data_0_8;
    assign token_in_vec_8[0] = token_0_8;
    assign in_chan_dep_vld_vec_8[1] = dep_chan_vld_1_8;
    assign in_chan_dep_data_vec_8[79 : 40] = dep_chan_data_1_8;
    assign token_in_vec_8[1] = token_1_8;
    assign in_chan_dep_vld_vec_8[2] = dep_chan_vld_3_8;
    assign in_chan_dep_data_vec_8[119 : 80] = dep_chan_data_3_8;
    assign token_in_vec_8[2] = token_3_8;
    assign in_chan_dep_vld_vec_8[3] = dep_chan_vld_6_8;
    assign in_chan_dep_data_vec_8[159 : 120] = dep_chan_data_6_8;
    assign token_in_vec_8[3] = token_6_8;
    assign in_chan_dep_vld_vec_8[4] = dep_chan_vld_7_8;
    assign in_chan_dep_data_vec_8[199 : 160] = dep_chan_data_7_8;
    assign token_in_vec_8[4] = token_7_8;
    assign in_chan_dep_vld_vec_8[5] = dep_chan_vld_9_8;
    assign in_chan_dep_data_vec_8[239 : 200] = dep_chan_data_9_8;
    assign token_in_vec_8[5] = token_9_8;
    assign in_chan_dep_vld_vec_8[6] = dep_chan_vld_10_8;
    assign in_chan_dep_data_vec_8[279 : 240] = dep_chan_data_10_8;
    assign token_in_vec_8[6] = token_10_8;
    assign in_chan_dep_vld_vec_8[7] = dep_chan_vld_11_8;
    assign in_chan_dep_data_vec_8[319 : 280] = dep_chan_data_11_8;
    assign token_in_vec_8[7] = token_11_8;
    assign in_chan_dep_vld_vec_8[8] = dep_chan_vld_12_8;
    assign in_chan_dep_data_vec_8[359 : 320] = dep_chan_data_12_8;
    assign token_in_vec_8[8] = token_12_8;
    assign in_chan_dep_vld_vec_8[9] = dep_chan_vld_13_8;
    assign in_chan_dep_data_vec_8[399 : 360] = dep_chan_data_13_8;
    assign token_in_vec_8[9] = token_13_8;
    assign in_chan_dep_vld_vec_8[10] = dep_chan_vld_14_8;
    assign in_chan_dep_data_vec_8[439 : 400] = dep_chan_data_14_8;
    assign token_in_vec_8[10] = token_14_8;
    assign in_chan_dep_vld_vec_8[11] = dep_chan_vld_15_8;
    assign in_chan_dep_data_vec_8[479 : 440] = dep_chan_data_15_8;
    assign token_in_vec_8[11] = token_15_8;
    assign in_chan_dep_vld_vec_8[12] = dep_chan_vld_16_8;
    assign in_chan_dep_data_vec_8[519 : 480] = dep_chan_data_16_8;
    assign token_in_vec_8[12] = token_16_8;
    assign in_chan_dep_vld_vec_8[13] = dep_chan_vld_17_8;
    assign in_chan_dep_data_vec_8[559 : 520] = dep_chan_data_17_8;
    assign token_in_vec_8[13] = token_17_8;
    assign in_chan_dep_vld_vec_8[14] = dep_chan_vld_18_8;
    assign in_chan_dep_data_vec_8[599 : 560] = dep_chan_data_18_8;
    assign token_in_vec_8[14] = token_18_8;
    assign in_chan_dep_vld_vec_8[15] = dep_chan_vld_19_8;
    assign in_chan_dep_data_vec_8[639 : 600] = dep_chan_data_19_8;
    assign token_in_vec_8[15] = token_19_8;
    assign in_chan_dep_vld_vec_8[16] = dep_chan_vld_20_8;
    assign in_chan_dep_data_vec_8[679 : 640] = dep_chan_data_20_8;
    assign token_in_vec_8[16] = token_20_8;
    assign in_chan_dep_vld_vec_8[17] = dep_chan_vld_21_8;
    assign in_chan_dep_data_vec_8[719 : 680] = dep_chan_data_21_8;
    assign token_in_vec_8[17] = token_21_8;
    assign in_chan_dep_vld_vec_8[18] = dep_chan_vld_22_8;
    assign in_chan_dep_data_vec_8[759 : 720] = dep_chan_data_22_8;
    assign token_in_vec_8[18] = token_22_8;
    assign in_chan_dep_vld_vec_8[19] = dep_chan_vld_23_8;
    assign in_chan_dep_data_vec_8[799 : 760] = dep_chan_data_23_8;
    assign token_in_vec_8[19] = token_23_8;
    assign in_chan_dep_vld_vec_8[20] = dep_chan_vld_24_8;
    assign in_chan_dep_data_vec_8[839 : 800] = dep_chan_data_24_8;
    assign token_in_vec_8[20] = token_24_8;
    assign in_chan_dep_vld_vec_8[21] = dep_chan_vld_25_8;
    assign in_chan_dep_data_vec_8[879 : 840] = dep_chan_data_25_8;
    assign token_in_vec_8[21] = token_25_8;
    assign in_chan_dep_vld_vec_8[22] = dep_chan_vld_26_8;
    assign in_chan_dep_data_vec_8[919 : 880] = dep_chan_data_26_8;
    assign token_in_vec_8[22] = token_26_8;
    assign in_chan_dep_vld_vec_8[23] = dep_chan_vld_27_8;
    assign in_chan_dep_data_vec_8[959 : 920] = dep_chan_data_27_8;
    assign token_in_vec_8[23] = token_27_8;
    assign in_chan_dep_vld_vec_8[24] = dep_chan_vld_28_8;
    assign in_chan_dep_data_vec_8[999 : 960] = dep_chan_data_28_8;
    assign token_in_vec_8[24] = token_28_8;
    assign in_chan_dep_vld_vec_8[25] = dep_chan_vld_29_8;
    assign in_chan_dep_data_vec_8[1039 : 1000] = dep_chan_data_29_8;
    assign token_in_vec_8[25] = token_29_8;
    assign in_chan_dep_vld_vec_8[26] = dep_chan_vld_30_8;
    assign in_chan_dep_data_vec_8[1079 : 1040] = dep_chan_data_30_8;
    assign token_in_vec_8[26] = token_30_8;
    assign in_chan_dep_vld_vec_8[27] = dep_chan_vld_31_8;
    assign in_chan_dep_data_vec_8[1119 : 1080] = dep_chan_data_31_8;
    assign token_in_vec_8[27] = token_31_8;
    assign in_chan_dep_vld_vec_8[28] = dep_chan_vld_32_8;
    assign in_chan_dep_data_vec_8[1159 : 1120] = dep_chan_data_32_8;
    assign token_in_vec_8[28] = token_32_8;
    assign in_chan_dep_vld_vec_8[29] = dep_chan_vld_33_8;
    assign in_chan_dep_data_vec_8[1199 : 1160] = dep_chan_data_33_8;
    assign token_in_vec_8[29] = token_33_8;
    assign in_chan_dep_vld_vec_8[30] = dep_chan_vld_34_8;
    assign in_chan_dep_data_vec_8[1239 : 1200] = dep_chan_data_34_8;
    assign token_in_vec_8[30] = token_34_8;
    assign in_chan_dep_vld_vec_8[31] = dep_chan_vld_35_8;
    assign in_chan_dep_data_vec_8[1279 : 1240] = dep_chan_data_35_8;
    assign token_in_vec_8[31] = token_35_8;
    assign in_chan_dep_vld_vec_8[32] = dep_chan_vld_36_8;
    assign in_chan_dep_data_vec_8[1319 : 1280] = dep_chan_data_36_8;
    assign token_in_vec_8[32] = token_36_8;
    assign dep_chan_vld_8_7 = out_chan_dep_vld_vec_8[0];
    assign dep_chan_data_8_7 = out_chan_dep_data_8;
    assign token_8_7 = token_out_vec_8[0];
    assign dep_chan_vld_8_9 = out_chan_dep_vld_vec_8[1];
    assign dep_chan_data_8_9 = out_chan_dep_data_8;
    assign token_8_9 = token_out_vec_8[1];
    assign dep_chan_vld_8_0 = out_chan_dep_vld_vec_8[2];
    assign dep_chan_data_8_0 = out_chan_dep_data_8;
    assign token_8_0 = token_out_vec_8[2];
    assign dep_chan_vld_8_1 = out_chan_dep_vld_vec_8[3];
    assign dep_chan_data_8_1 = out_chan_dep_data_8;
    assign token_8_1 = token_out_vec_8[3];
    assign dep_chan_vld_8_3 = out_chan_dep_vld_vec_8[4];
    assign dep_chan_data_8_3 = out_chan_dep_data_8;
    assign token_8_3 = token_out_vec_8[4];
    assign dep_chan_vld_8_6 = out_chan_dep_vld_vec_8[5];
    assign dep_chan_data_8_6 = out_chan_dep_data_8;
    assign token_8_6 = token_out_vec_8[5];
    assign dep_chan_vld_8_10 = out_chan_dep_vld_vec_8[6];
    assign dep_chan_data_8_10 = out_chan_dep_data_8;
    assign token_8_10 = token_out_vec_8[6];
    assign dep_chan_vld_8_11 = out_chan_dep_vld_vec_8[7];
    assign dep_chan_data_8_11 = out_chan_dep_data_8;
    assign token_8_11 = token_out_vec_8[7];
    assign dep_chan_vld_8_12 = out_chan_dep_vld_vec_8[8];
    assign dep_chan_data_8_12 = out_chan_dep_data_8;
    assign token_8_12 = token_out_vec_8[8];
    assign dep_chan_vld_8_13 = out_chan_dep_vld_vec_8[9];
    assign dep_chan_data_8_13 = out_chan_dep_data_8;
    assign token_8_13 = token_out_vec_8[9];
    assign dep_chan_vld_8_14 = out_chan_dep_vld_vec_8[10];
    assign dep_chan_data_8_14 = out_chan_dep_data_8;
    assign token_8_14 = token_out_vec_8[10];
    assign dep_chan_vld_8_15 = out_chan_dep_vld_vec_8[11];
    assign dep_chan_data_8_15 = out_chan_dep_data_8;
    assign token_8_15 = token_out_vec_8[11];
    assign dep_chan_vld_8_16 = out_chan_dep_vld_vec_8[12];
    assign dep_chan_data_8_16 = out_chan_dep_data_8;
    assign token_8_16 = token_out_vec_8[12];
    assign dep_chan_vld_8_17 = out_chan_dep_vld_vec_8[13];
    assign dep_chan_data_8_17 = out_chan_dep_data_8;
    assign token_8_17 = token_out_vec_8[13];
    assign dep_chan_vld_8_18 = out_chan_dep_vld_vec_8[14];
    assign dep_chan_data_8_18 = out_chan_dep_data_8;
    assign token_8_18 = token_out_vec_8[14];
    assign dep_chan_vld_8_19 = out_chan_dep_vld_vec_8[15];
    assign dep_chan_data_8_19 = out_chan_dep_data_8;
    assign token_8_19 = token_out_vec_8[15];
    assign dep_chan_vld_8_20 = out_chan_dep_vld_vec_8[16];
    assign dep_chan_data_8_20 = out_chan_dep_data_8;
    assign token_8_20 = token_out_vec_8[16];
    assign dep_chan_vld_8_21 = out_chan_dep_vld_vec_8[17];
    assign dep_chan_data_8_21 = out_chan_dep_data_8;
    assign token_8_21 = token_out_vec_8[17];
    assign dep_chan_vld_8_22 = out_chan_dep_vld_vec_8[18];
    assign dep_chan_data_8_22 = out_chan_dep_data_8;
    assign token_8_22 = token_out_vec_8[18];
    assign dep_chan_vld_8_23 = out_chan_dep_vld_vec_8[19];
    assign dep_chan_data_8_23 = out_chan_dep_data_8;
    assign token_8_23 = token_out_vec_8[19];
    assign dep_chan_vld_8_24 = out_chan_dep_vld_vec_8[20];
    assign dep_chan_data_8_24 = out_chan_dep_data_8;
    assign token_8_24 = token_out_vec_8[20];
    assign dep_chan_vld_8_25 = out_chan_dep_vld_vec_8[21];
    assign dep_chan_data_8_25 = out_chan_dep_data_8;
    assign token_8_25 = token_out_vec_8[21];
    assign dep_chan_vld_8_26 = out_chan_dep_vld_vec_8[22];
    assign dep_chan_data_8_26 = out_chan_dep_data_8;
    assign token_8_26 = token_out_vec_8[22];
    assign dep_chan_vld_8_27 = out_chan_dep_vld_vec_8[23];
    assign dep_chan_data_8_27 = out_chan_dep_data_8;
    assign token_8_27 = token_out_vec_8[23];
    assign dep_chan_vld_8_28 = out_chan_dep_vld_vec_8[24];
    assign dep_chan_data_8_28 = out_chan_dep_data_8;
    assign token_8_28 = token_out_vec_8[24];
    assign dep_chan_vld_8_29 = out_chan_dep_vld_vec_8[25];
    assign dep_chan_data_8_29 = out_chan_dep_data_8;
    assign token_8_29 = token_out_vec_8[25];
    assign dep_chan_vld_8_30 = out_chan_dep_vld_vec_8[26];
    assign dep_chan_data_8_30 = out_chan_dep_data_8;
    assign token_8_30 = token_out_vec_8[26];
    assign dep_chan_vld_8_31 = out_chan_dep_vld_vec_8[27];
    assign dep_chan_data_8_31 = out_chan_dep_data_8;
    assign token_8_31 = token_out_vec_8[27];
    assign dep_chan_vld_8_32 = out_chan_dep_vld_vec_8[28];
    assign dep_chan_data_8_32 = out_chan_dep_data_8;
    assign token_8_32 = token_out_vec_8[28];
    assign dep_chan_vld_8_33 = out_chan_dep_vld_vec_8[29];
    assign dep_chan_data_8_33 = out_chan_dep_data_8;
    assign token_8_33 = token_out_vec_8[29];
    assign dep_chan_vld_8_34 = out_chan_dep_vld_vec_8[30];
    assign dep_chan_data_8_34 = out_chan_dep_data_8;
    assign token_8_34 = token_out_vec_8[30];
    assign dep_chan_vld_8_35 = out_chan_dep_vld_vec_8[31];
    assign dep_chan_data_8_35 = out_chan_dep_data_8;
    assign token_8_35 = token_out_vec_8[31];
    assign dep_chan_vld_8_36 = out_chan_dep_vld_vec_8[32];
    assign dep_chan_data_8_36 = out_chan_dep_data_8;
    assign token_8_36 = token_out_vec_8[32];

    // Process: ProcessingElement_4_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 9, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_9 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_9),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_9),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_9),
        .token_in_vec(token_in_vec_9),
        .dl_detect_in(dl_detect_out),
        .origin(origin[9]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_9),
        .out_chan_dep_data(out_chan_dep_data_9),
        .token_out_vec(token_out_vec_9),
        .dl_detect_out(dl_in_vec[9]));

    assign proc_9_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_3_blk_n) | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_3_blk_n) | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_WriteC_Flattened_fu_179.cPipes_3_blk_n);
    assign proc_9_data_PIPO_blk[0] = 1'b0;
    assign proc_9_start_FIFO_blk[0] = 1'b0;
    assign proc_9_TLF_FIFO_blk[0] = 1'b0;
    assign proc_9_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_9_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_9[0] = dl_detect_out ? proc_dep_vld_vec_9_reg[0] : (proc_9_data_FIFO_blk[0] | proc_9_data_PIPO_blk[0] | proc_9_start_FIFO_blk[0] | proc_9_TLF_FIFO_blk[0] | proc_9_input_sync_blk[0] | proc_9_output_sync_blk[0]);
    assign proc_9_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_4_blk_n) | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_4_blk_n) | (~ProcessingElement_4_U0.grp_ProcessingElement_4_Pipeline_WriteC_Flattened_fu_179.cPipes_4_blk_n);
    assign proc_9_data_PIPO_blk[1] = 1'b0;
    assign proc_9_start_FIFO_blk[1] = 1'b0;
    assign proc_9_TLF_FIFO_blk[1] = 1'b0;
    assign proc_9_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_9_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_9[1] = dl_detect_out ? proc_dep_vld_vec_9_reg[1] : (proc_9_data_FIFO_blk[1] | proc_9_data_PIPO_blk[1] | proc_9_start_FIFO_blk[1] | proc_9_TLF_FIFO_blk[1] | proc_9_input_sync_blk[1] | proc_9_output_sync_blk[1]);
    assign proc_9_data_FIFO_blk[2] = 1'b0;
    assign proc_9_data_PIPO_blk[2] = 1'b0;
    assign proc_9_start_FIFO_blk[2] = 1'b0;
    assign proc_9_TLF_FIFO_blk[2] = 1'b0;
    assign proc_9_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_9_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_9[2] = dl_detect_out ? proc_dep_vld_vec_9_reg[2] : (proc_9_data_FIFO_blk[2] | proc_9_data_PIPO_blk[2] | proc_9_start_FIFO_blk[2] | proc_9_TLF_FIFO_blk[2] | proc_9_input_sync_blk[2] | proc_9_output_sync_blk[2]);
    assign proc_9_data_FIFO_blk[3] = 1'b0;
    assign proc_9_data_PIPO_blk[3] = 1'b0;
    assign proc_9_start_FIFO_blk[3] = 1'b0;
    assign proc_9_TLF_FIFO_blk[3] = 1'b0;
    assign proc_9_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_9_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_9[3] = dl_detect_out ? proc_dep_vld_vec_9_reg[3] : (proc_9_data_FIFO_blk[3] | proc_9_data_PIPO_blk[3] | proc_9_start_FIFO_blk[3] | proc_9_TLF_FIFO_blk[3] | proc_9_input_sync_blk[3] | proc_9_output_sync_blk[3]);
    assign proc_9_data_FIFO_blk[4] = 1'b0;
    assign proc_9_data_PIPO_blk[4] = 1'b0;
    assign proc_9_start_FIFO_blk[4] = 1'b0;
    assign proc_9_TLF_FIFO_blk[4] = 1'b0;
    assign proc_9_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_9_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_9[4] = dl_detect_out ? proc_dep_vld_vec_9_reg[4] : (proc_9_data_FIFO_blk[4] | proc_9_data_PIPO_blk[4] | proc_9_start_FIFO_blk[4] | proc_9_TLF_FIFO_blk[4] | proc_9_input_sync_blk[4] | proc_9_output_sync_blk[4]);
    assign proc_9_data_FIFO_blk[5] = 1'b0;
    assign proc_9_data_PIPO_blk[5] = 1'b0;
    assign proc_9_start_FIFO_blk[5] = 1'b0;
    assign proc_9_TLF_FIFO_blk[5] = 1'b0;
    assign proc_9_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_9_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_9[5] = dl_detect_out ? proc_dep_vld_vec_9_reg[5] : (proc_9_data_FIFO_blk[5] | proc_9_data_PIPO_blk[5] | proc_9_start_FIFO_blk[5] | proc_9_TLF_FIFO_blk[5] | proc_9_input_sync_blk[5] | proc_9_output_sync_blk[5]);
    assign proc_9_data_FIFO_blk[6] = 1'b0;
    assign proc_9_data_PIPO_blk[6] = 1'b0;
    assign proc_9_start_FIFO_blk[6] = 1'b0;
    assign proc_9_TLF_FIFO_blk[6] = 1'b0;
    assign proc_9_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_9_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_9[6] = dl_detect_out ? proc_dep_vld_vec_9_reg[6] : (proc_9_data_FIFO_blk[6] | proc_9_data_PIPO_blk[6] | proc_9_start_FIFO_blk[6] | proc_9_TLF_FIFO_blk[6] | proc_9_input_sync_blk[6] | proc_9_output_sync_blk[6]);
    assign proc_9_data_FIFO_blk[7] = 1'b0;
    assign proc_9_data_PIPO_blk[7] = 1'b0;
    assign proc_9_start_FIFO_blk[7] = 1'b0;
    assign proc_9_TLF_FIFO_blk[7] = 1'b0;
    assign proc_9_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_9_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_9[7] = dl_detect_out ? proc_dep_vld_vec_9_reg[7] : (proc_9_data_FIFO_blk[7] | proc_9_data_PIPO_blk[7] | proc_9_start_FIFO_blk[7] | proc_9_TLF_FIFO_blk[7] | proc_9_input_sync_blk[7] | proc_9_output_sync_blk[7]);
    assign proc_9_data_FIFO_blk[8] = 1'b0;
    assign proc_9_data_PIPO_blk[8] = 1'b0;
    assign proc_9_start_FIFO_blk[8] = 1'b0;
    assign proc_9_TLF_FIFO_blk[8] = 1'b0;
    assign proc_9_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_9_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_9[8] = dl_detect_out ? proc_dep_vld_vec_9_reg[8] : (proc_9_data_FIFO_blk[8] | proc_9_data_PIPO_blk[8] | proc_9_start_FIFO_blk[8] | proc_9_TLF_FIFO_blk[8] | proc_9_input_sync_blk[8] | proc_9_output_sync_blk[8]);
    assign proc_9_data_FIFO_blk[9] = 1'b0;
    assign proc_9_data_PIPO_blk[9] = 1'b0;
    assign proc_9_start_FIFO_blk[9] = 1'b0;
    assign proc_9_TLF_FIFO_blk[9] = 1'b0;
    assign proc_9_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_9_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_9[9] = dl_detect_out ? proc_dep_vld_vec_9_reg[9] : (proc_9_data_FIFO_blk[9] | proc_9_data_PIPO_blk[9] | proc_9_start_FIFO_blk[9] | proc_9_TLF_FIFO_blk[9] | proc_9_input_sync_blk[9] | proc_9_output_sync_blk[9]);
    assign proc_9_data_FIFO_blk[10] = 1'b0;
    assign proc_9_data_PIPO_blk[10] = 1'b0;
    assign proc_9_start_FIFO_blk[10] = 1'b0;
    assign proc_9_TLF_FIFO_blk[10] = 1'b0;
    assign proc_9_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_9_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_9[10] = dl_detect_out ? proc_dep_vld_vec_9_reg[10] : (proc_9_data_FIFO_blk[10] | proc_9_data_PIPO_blk[10] | proc_9_start_FIFO_blk[10] | proc_9_TLF_FIFO_blk[10] | proc_9_input_sync_blk[10] | proc_9_output_sync_blk[10]);
    assign proc_9_data_FIFO_blk[11] = 1'b0;
    assign proc_9_data_PIPO_blk[11] = 1'b0;
    assign proc_9_start_FIFO_blk[11] = 1'b0;
    assign proc_9_TLF_FIFO_blk[11] = 1'b0;
    assign proc_9_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_9_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_9[11] = dl_detect_out ? proc_dep_vld_vec_9_reg[11] : (proc_9_data_FIFO_blk[11] | proc_9_data_PIPO_blk[11] | proc_9_start_FIFO_blk[11] | proc_9_TLF_FIFO_blk[11] | proc_9_input_sync_blk[11] | proc_9_output_sync_blk[11]);
    assign proc_9_data_FIFO_blk[12] = 1'b0;
    assign proc_9_data_PIPO_blk[12] = 1'b0;
    assign proc_9_start_FIFO_blk[12] = 1'b0;
    assign proc_9_TLF_FIFO_blk[12] = 1'b0;
    assign proc_9_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_9_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_9[12] = dl_detect_out ? proc_dep_vld_vec_9_reg[12] : (proc_9_data_FIFO_blk[12] | proc_9_data_PIPO_blk[12] | proc_9_start_FIFO_blk[12] | proc_9_TLF_FIFO_blk[12] | proc_9_input_sync_blk[12] | proc_9_output_sync_blk[12]);
    assign proc_9_data_FIFO_blk[13] = 1'b0;
    assign proc_9_data_PIPO_blk[13] = 1'b0;
    assign proc_9_start_FIFO_blk[13] = 1'b0;
    assign proc_9_TLF_FIFO_blk[13] = 1'b0;
    assign proc_9_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_9_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_9[13] = dl_detect_out ? proc_dep_vld_vec_9_reg[13] : (proc_9_data_FIFO_blk[13] | proc_9_data_PIPO_blk[13] | proc_9_start_FIFO_blk[13] | proc_9_TLF_FIFO_blk[13] | proc_9_input_sync_blk[13] | proc_9_output_sync_blk[13]);
    assign proc_9_data_FIFO_blk[14] = 1'b0;
    assign proc_9_data_PIPO_blk[14] = 1'b0;
    assign proc_9_start_FIFO_blk[14] = 1'b0;
    assign proc_9_TLF_FIFO_blk[14] = 1'b0;
    assign proc_9_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_9_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_9[14] = dl_detect_out ? proc_dep_vld_vec_9_reg[14] : (proc_9_data_FIFO_blk[14] | proc_9_data_PIPO_blk[14] | proc_9_start_FIFO_blk[14] | proc_9_TLF_FIFO_blk[14] | proc_9_input_sync_blk[14] | proc_9_output_sync_blk[14]);
    assign proc_9_data_FIFO_blk[15] = 1'b0;
    assign proc_9_data_PIPO_blk[15] = 1'b0;
    assign proc_9_start_FIFO_blk[15] = 1'b0;
    assign proc_9_TLF_FIFO_blk[15] = 1'b0;
    assign proc_9_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_9_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_9[15] = dl_detect_out ? proc_dep_vld_vec_9_reg[15] : (proc_9_data_FIFO_blk[15] | proc_9_data_PIPO_blk[15] | proc_9_start_FIFO_blk[15] | proc_9_TLF_FIFO_blk[15] | proc_9_input_sync_blk[15] | proc_9_output_sync_blk[15]);
    assign proc_9_data_FIFO_blk[16] = 1'b0;
    assign proc_9_data_PIPO_blk[16] = 1'b0;
    assign proc_9_start_FIFO_blk[16] = 1'b0;
    assign proc_9_TLF_FIFO_blk[16] = 1'b0;
    assign proc_9_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_9_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_9[16] = dl_detect_out ? proc_dep_vld_vec_9_reg[16] : (proc_9_data_FIFO_blk[16] | proc_9_data_PIPO_blk[16] | proc_9_start_FIFO_blk[16] | proc_9_TLF_FIFO_blk[16] | proc_9_input_sync_blk[16] | proc_9_output_sync_blk[16]);
    assign proc_9_data_FIFO_blk[17] = 1'b0;
    assign proc_9_data_PIPO_blk[17] = 1'b0;
    assign proc_9_start_FIFO_blk[17] = 1'b0;
    assign proc_9_TLF_FIFO_blk[17] = 1'b0;
    assign proc_9_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_9_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_9[17] = dl_detect_out ? proc_dep_vld_vec_9_reg[17] : (proc_9_data_FIFO_blk[17] | proc_9_data_PIPO_blk[17] | proc_9_start_FIFO_blk[17] | proc_9_TLF_FIFO_blk[17] | proc_9_input_sync_blk[17] | proc_9_output_sync_blk[17]);
    assign proc_9_data_FIFO_blk[18] = 1'b0;
    assign proc_9_data_PIPO_blk[18] = 1'b0;
    assign proc_9_start_FIFO_blk[18] = 1'b0;
    assign proc_9_TLF_FIFO_blk[18] = 1'b0;
    assign proc_9_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_9_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_9[18] = dl_detect_out ? proc_dep_vld_vec_9_reg[18] : (proc_9_data_FIFO_blk[18] | proc_9_data_PIPO_blk[18] | proc_9_start_FIFO_blk[18] | proc_9_TLF_FIFO_blk[18] | proc_9_input_sync_blk[18] | proc_9_output_sync_blk[18]);
    assign proc_9_data_FIFO_blk[19] = 1'b0;
    assign proc_9_data_PIPO_blk[19] = 1'b0;
    assign proc_9_start_FIFO_blk[19] = 1'b0;
    assign proc_9_TLF_FIFO_blk[19] = 1'b0;
    assign proc_9_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_9_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_9[19] = dl_detect_out ? proc_dep_vld_vec_9_reg[19] : (proc_9_data_FIFO_blk[19] | proc_9_data_PIPO_blk[19] | proc_9_start_FIFO_blk[19] | proc_9_TLF_FIFO_blk[19] | proc_9_input_sync_blk[19] | proc_9_output_sync_blk[19]);
    assign proc_9_data_FIFO_blk[20] = 1'b0;
    assign proc_9_data_PIPO_blk[20] = 1'b0;
    assign proc_9_start_FIFO_blk[20] = 1'b0;
    assign proc_9_TLF_FIFO_blk[20] = 1'b0;
    assign proc_9_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_9_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_9[20] = dl_detect_out ? proc_dep_vld_vec_9_reg[20] : (proc_9_data_FIFO_blk[20] | proc_9_data_PIPO_blk[20] | proc_9_start_FIFO_blk[20] | proc_9_TLF_FIFO_blk[20] | proc_9_input_sync_blk[20] | proc_9_output_sync_blk[20]);
    assign proc_9_data_FIFO_blk[21] = 1'b0;
    assign proc_9_data_PIPO_blk[21] = 1'b0;
    assign proc_9_start_FIFO_blk[21] = 1'b0;
    assign proc_9_TLF_FIFO_blk[21] = 1'b0;
    assign proc_9_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_9_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_9[21] = dl_detect_out ? proc_dep_vld_vec_9_reg[21] : (proc_9_data_FIFO_blk[21] | proc_9_data_PIPO_blk[21] | proc_9_start_FIFO_blk[21] | proc_9_TLF_FIFO_blk[21] | proc_9_input_sync_blk[21] | proc_9_output_sync_blk[21]);
    assign proc_9_data_FIFO_blk[22] = 1'b0;
    assign proc_9_data_PIPO_blk[22] = 1'b0;
    assign proc_9_start_FIFO_blk[22] = 1'b0;
    assign proc_9_TLF_FIFO_blk[22] = 1'b0;
    assign proc_9_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_9_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_9[22] = dl_detect_out ? proc_dep_vld_vec_9_reg[22] : (proc_9_data_FIFO_blk[22] | proc_9_data_PIPO_blk[22] | proc_9_start_FIFO_blk[22] | proc_9_TLF_FIFO_blk[22] | proc_9_input_sync_blk[22] | proc_9_output_sync_blk[22]);
    assign proc_9_data_FIFO_blk[23] = 1'b0;
    assign proc_9_data_PIPO_blk[23] = 1'b0;
    assign proc_9_start_FIFO_blk[23] = 1'b0;
    assign proc_9_TLF_FIFO_blk[23] = 1'b0;
    assign proc_9_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_9_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_9[23] = dl_detect_out ? proc_dep_vld_vec_9_reg[23] : (proc_9_data_FIFO_blk[23] | proc_9_data_PIPO_blk[23] | proc_9_start_FIFO_blk[23] | proc_9_TLF_FIFO_blk[23] | proc_9_input_sync_blk[23] | proc_9_output_sync_blk[23]);
    assign proc_9_data_FIFO_blk[24] = 1'b0;
    assign proc_9_data_PIPO_blk[24] = 1'b0;
    assign proc_9_start_FIFO_blk[24] = 1'b0;
    assign proc_9_TLF_FIFO_blk[24] = 1'b0;
    assign proc_9_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_9_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_9[24] = dl_detect_out ? proc_dep_vld_vec_9_reg[24] : (proc_9_data_FIFO_blk[24] | proc_9_data_PIPO_blk[24] | proc_9_start_FIFO_blk[24] | proc_9_TLF_FIFO_blk[24] | proc_9_input_sync_blk[24] | proc_9_output_sync_blk[24]);
    assign proc_9_data_FIFO_blk[25] = 1'b0;
    assign proc_9_data_PIPO_blk[25] = 1'b0;
    assign proc_9_start_FIFO_blk[25] = 1'b0;
    assign proc_9_TLF_FIFO_blk[25] = 1'b0;
    assign proc_9_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_9_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_9[25] = dl_detect_out ? proc_dep_vld_vec_9_reg[25] : (proc_9_data_FIFO_blk[25] | proc_9_data_PIPO_blk[25] | proc_9_start_FIFO_blk[25] | proc_9_TLF_FIFO_blk[25] | proc_9_input_sync_blk[25] | proc_9_output_sync_blk[25]);
    assign proc_9_data_FIFO_blk[26] = 1'b0;
    assign proc_9_data_PIPO_blk[26] = 1'b0;
    assign proc_9_start_FIFO_blk[26] = 1'b0;
    assign proc_9_TLF_FIFO_blk[26] = 1'b0;
    assign proc_9_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_9_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_9[26] = dl_detect_out ? proc_dep_vld_vec_9_reg[26] : (proc_9_data_FIFO_blk[26] | proc_9_data_PIPO_blk[26] | proc_9_start_FIFO_blk[26] | proc_9_TLF_FIFO_blk[26] | proc_9_input_sync_blk[26] | proc_9_output_sync_blk[26]);
    assign proc_9_data_FIFO_blk[27] = 1'b0;
    assign proc_9_data_PIPO_blk[27] = 1'b0;
    assign proc_9_start_FIFO_blk[27] = 1'b0;
    assign proc_9_TLF_FIFO_blk[27] = 1'b0;
    assign proc_9_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_9_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_9[27] = dl_detect_out ? proc_dep_vld_vec_9_reg[27] : (proc_9_data_FIFO_blk[27] | proc_9_data_PIPO_blk[27] | proc_9_start_FIFO_blk[27] | proc_9_TLF_FIFO_blk[27] | proc_9_input_sync_blk[27] | proc_9_output_sync_blk[27]);
    assign proc_9_data_FIFO_blk[28] = 1'b0;
    assign proc_9_data_PIPO_blk[28] = 1'b0;
    assign proc_9_start_FIFO_blk[28] = 1'b0;
    assign proc_9_TLF_FIFO_blk[28] = 1'b0;
    assign proc_9_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_9_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_9[28] = dl_detect_out ? proc_dep_vld_vec_9_reg[28] : (proc_9_data_FIFO_blk[28] | proc_9_data_PIPO_blk[28] | proc_9_start_FIFO_blk[28] | proc_9_TLF_FIFO_blk[28] | proc_9_input_sync_blk[28] | proc_9_output_sync_blk[28]);
    assign proc_9_data_FIFO_blk[29] = 1'b0;
    assign proc_9_data_PIPO_blk[29] = 1'b0;
    assign proc_9_start_FIFO_blk[29] = 1'b0;
    assign proc_9_TLF_FIFO_blk[29] = 1'b0;
    assign proc_9_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_9_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_9[29] = dl_detect_out ? proc_dep_vld_vec_9_reg[29] : (proc_9_data_FIFO_blk[29] | proc_9_data_PIPO_blk[29] | proc_9_start_FIFO_blk[29] | proc_9_TLF_FIFO_blk[29] | proc_9_input_sync_blk[29] | proc_9_output_sync_blk[29]);
    assign proc_9_data_FIFO_blk[30] = 1'b0;
    assign proc_9_data_PIPO_blk[30] = 1'b0;
    assign proc_9_start_FIFO_blk[30] = 1'b0;
    assign proc_9_TLF_FIFO_blk[30] = 1'b0;
    assign proc_9_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_9_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_9[30] = dl_detect_out ? proc_dep_vld_vec_9_reg[30] : (proc_9_data_FIFO_blk[30] | proc_9_data_PIPO_blk[30] | proc_9_start_FIFO_blk[30] | proc_9_TLF_FIFO_blk[30] | proc_9_input_sync_blk[30] | proc_9_output_sync_blk[30]);
    assign proc_9_data_FIFO_blk[31] = 1'b0;
    assign proc_9_data_PIPO_blk[31] = 1'b0;
    assign proc_9_start_FIFO_blk[31] = 1'b0;
    assign proc_9_TLF_FIFO_blk[31] = 1'b0;
    assign proc_9_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_9_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_9[31] = dl_detect_out ? proc_dep_vld_vec_9_reg[31] : (proc_9_data_FIFO_blk[31] | proc_9_data_PIPO_blk[31] | proc_9_start_FIFO_blk[31] | proc_9_TLF_FIFO_blk[31] | proc_9_input_sync_blk[31] | proc_9_output_sync_blk[31]);
    assign proc_9_data_FIFO_blk[32] = 1'b0;
    assign proc_9_data_PIPO_blk[32] = 1'b0;
    assign proc_9_start_FIFO_blk[32] = 1'b0;
    assign proc_9_TLF_FIFO_blk[32] = 1'b0;
    assign proc_9_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_4_U0_ap_ready & ProcessingElement_4_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_9_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_9[32] = dl_detect_out ? proc_dep_vld_vec_9_reg[32] : (proc_9_data_FIFO_blk[32] | proc_9_data_PIPO_blk[32] | proc_9_start_FIFO_blk[32] | proc_9_TLF_FIFO_blk[32] | proc_9_input_sync_blk[32] | proc_9_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_9_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_9_reg <= proc_dep_vld_vec_9;
        end
    end
    assign in_chan_dep_vld_vec_9[0] = dep_chan_vld_0_9;
    assign in_chan_dep_data_vec_9[39 : 0] = dep_chan_data_0_9;
    assign token_in_vec_9[0] = token_0_9;
    assign in_chan_dep_vld_vec_9[1] = dep_chan_vld_1_9;
    assign in_chan_dep_data_vec_9[79 : 40] = dep_chan_data_1_9;
    assign token_in_vec_9[1] = token_1_9;
    assign in_chan_dep_vld_vec_9[2] = dep_chan_vld_3_9;
    assign in_chan_dep_data_vec_9[119 : 80] = dep_chan_data_3_9;
    assign token_in_vec_9[2] = token_3_9;
    assign in_chan_dep_vld_vec_9[3] = dep_chan_vld_6_9;
    assign in_chan_dep_data_vec_9[159 : 120] = dep_chan_data_6_9;
    assign token_in_vec_9[3] = token_6_9;
    assign in_chan_dep_vld_vec_9[4] = dep_chan_vld_7_9;
    assign in_chan_dep_data_vec_9[199 : 160] = dep_chan_data_7_9;
    assign token_in_vec_9[4] = token_7_9;
    assign in_chan_dep_vld_vec_9[5] = dep_chan_vld_8_9;
    assign in_chan_dep_data_vec_9[239 : 200] = dep_chan_data_8_9;
    assign token_in_vec_9[5] = token_8_9;
    assign in_chan_dep_vld_vec_9[6] = dep_chan_vld_10_9;
    assign in_chan_dep_data_vec_9[279 : 240] = dep_chan_data_10_9;
    assign token_in_vec_9[6] = token_10_9;
    assign in_chan_dep_vld_vec_9[7] = dep_chan_vld_11_9;
    assign in_chan_dep_data_vec_9[319 : 280] = dep_chan_data_11_9;
    assign token_in_vec_9[7] = token_11_9;
    assign in_chan_dep_vld_vec_9[8] = dep_chan_vld_12_9;
    assign in_chan_dep_data_vec_9[359 : 320] = dep_chan_data_12_9;
    assign token_in_vec_9[8] = token_12_9;
    assign in_chan_dep_vld_vec_9[9] = dep_chan_vld_13_9;
    assign in_chan_dep_data_vec_9[399 : 360] = dep_chan_data_13_9;
    assign token_in_vec_9[9] = token_13_9;
    assign in_chan_dep_vld_vec_9[10] = dep_chan_vld_14_9;
    assign in_chan_dep_data_vec_9[439 : 400] = dep_chan_data_14_9;
    assign token_in_vec_9[10] = token_14_9;
    assign in_chan_dep_vld_vec_9[11] = dep_chan_vld_15_9;
    assign in_chan_dep_data_vec_9[479 : 440] = dep_chan_data_15_9;
    assign token_in_vec_9[11] = token_15_9;
    assign in_chan_dep_vld_vec_9[12] = dep_chan_vld_16_9;
    assign in_chan_dep_data_vec_9[519 : 480] = dep_chan_data_16_9;
    assign token_in_vec_9[12] = token_16_9;
    assign in_chan_dep_vld_vec_9[13] = dep_chan_vld_17_9;
    assign in_chan_dep_data_vec_9[559 : 520] = dep_chan_data_17_9;
    assign token_in_vec_9[13] = token_17_9;
    assign in_chan_dep_vld_vec_9[14] = dep_chan_vld_18_9;
    assign in_chan_dep_data_vec_9[599 : 560] = dep_chan_data_18_9;
    assign token_in_vec_9[14] = token_18_9;
    assign in_chan_dep_vld_vec_9[15] = dep_chan_vld_19_9;
    assign in_chan_dep_data_vec_9[639 : 600] = dep_chan_data_19_9;
    assign token_in_vec_9[15] = token_19_9;
    assign in_chan_dep_vld_vec_9[16] = dep_chan_vld_20_9;
    assign in_chan_dep_data_vec_9[679 : 640] = dep_chan_data_20_9;
    assign token_in_vec_9[16] = token_20_9;
    assign in_chan_dep_vld_vec_9[17] = dep_chan_vld_21_9;
    assign in_chan_dep_data_vec_9[719 : 680] = dep_chan_data_21_9;
    assign token_in_vec_9[17] = token_21_9;
    assign in_chan_dep_vld_vec_9[18] = dep_chan_vld_22_9;
    assign in_chan_dep_data_vec_9[759 : 720] = dep_chan_data_22_9;
    assign token_in_vec_9[18] = token_22_9;
    assign in_chan_dep_vld_vec_9[19] = dep_chan_vld_23_9;
    assign in_chan_dep_data_vec_9[799 : 760] = dep_chan_data_23_9;
    assign token_in_vec_9[19] = token_23_9;
    assign in_chan_dep_vld_vec_9[20] = dep_chan_vld_24_9;
    assign in_chan_dep_data_vec_9[839 : 800] = dep_chan_data_24_9;
    assign token_in_vec_9[20] = token_24_9;
    assign in_chan_dep_vld_vec_9[21] = dep_chan_vld_25_9;
    assign in_chan_dep_data_vec_9[879 : 840] = dep_chan_data_25_9;
    assign token_in_vec_9[21] = token_25_9;
    assign in_chan_dep_vld_vec_9[22] = dep_chan_vld_26_9;
    assign in_chan_dep_data_vec_9[919 : 880] = dep_chan_data_26_9;
    assign token_in_vec_9[22] = token_26_9;
    assign in_chan_dep_vld_vec_9[23] = dep_chan_vld_27_9;
    assign in_chan_dep_data_vec_9[959 : 920] = dep_chan_data_27_9;
    assign token_in_vec_9[23] = token_27_9;
    assign in_chan_dep_vld_vec_9[24] = dep_chan_vld_28_9;
    assign in_chan_dep_data_vec_9[999 : 960] = dep_chan_data_28_9;
    assign token_in_vec_9[24] = token_28_9;
    assign in_chan_dep_vld_vec_9[25] = dep_chan_vld_29_9;
    assign in_chan_dep_data_vec_9[1039 : 1000] = dep_chan_data_29_9;
    assign token_in_vec_9[25] = token_29_9;
    assign in_chan_dep_vld_vec_9[26] = dep_chan_vld_30_9;
    assign in_chan_dep_data_vec_9[1079 : 1040] = dep_chan_data_30_9;
    assign token_in_vec_9[26] = token_30_9;
    assign in_chan_dep_vld_vec_9[27] = dep_chan_vld_31_9;
    assign in_chan_dep_data_vec_9[1119 : 1080] = dep_chan_data_31_9;
    assign token_in_vec_9[27] = token_31_9;
    assign in_chan_dep_vld_vec_9[28] = dep_chan_vld_32_9;
    assign in_chan_dep_data_vec_9[1159 : 1120] = dep_chan_data_32_9;
    assign token_in_vec_9[28] = token_32_9;
    assign in_chan_dep_vld_vec_9[29] = dep_chan_vld_33_9;
    assign in_chan_dep_data_vec_9[1199 : 1160] = dep_chan_data_33_9;
    assign token_in_vec_9[29] = token_33_9;
    assign in_chan_dep_vld_vec_9[30] = dep_chan_vld_34_9;
    assign in_chan_dep_data_vec_9[1239 : 1200] = dep_chan_data_34_9;
    assign token_in_vec_9[30] = token_34_9;
    assign in_chan_dep_vld_vec_9[31] = dep_chan_vld_35_9;
    assign in_chan_dep_data_vec_9[1279 : 1240] = dep_chan_data_35_9;
    assign token_in_vec_9[31] = token_35_9;
    assign in_chan_dep_vld_vec_9[32] = dep_chan_vld_36_9;
    assign in_chan_dep_data_vec_9[1319 : 1280] = dep_chan_data_36_9;
    assign token_in_vec_9[32] = token_36_9;
    assign dep_chan_vld_9_8 = out_chan_dep_vld_vec_9[0];
    assign dep_chan_data_9_8 = out_chan_dep_data_9;
    assign token_9_8 = token_out_vec_9[0];
    assign dep_chan_vld_9_10 = out_chan_dep_vld_vec_9[1];
    assign dep_chan_data_9_10 = out_chan_dep_data_9;
    assign token_9_10 = token_out_vec_9[1];
    assign dep_chan_vld_9_0 = out_chan_dep_vld_vec_9[2];
    assign dep_chan_data_9_0 = out_chan_dep_data_9;
    assign token_9_0 = token_out_vec_9[2];
    assign dep_chan_vld_9_1 = out_chan_dep_vld_vec_9[3];
    assign dep_chan_data_9_1 = out_chan_dep_data_9;
    assign token_9_1 = token_out_vec_9[3];
    assign dep_chan_vld_9_3 = out_chan_dep_vld_vec_9[4];
    assign dep_chan_data_9_3 = out_chan_dep_data_9;
    assign token_9_3 = token_out_vec_9[4];
    assign dep_chan_vld_9_6 = out_chan_dep_vld_vec_9[5];
    assign dep_chan_data_9_6 = out_chan_dep_data_9;
    assign token_9_6 = token_out_vec_9[5];
    assign dep_chan_vld_9_7 = out_chan_dep_vld_vec_9[6];
    assign dep_chan_data_9_7 = out_chan_dep_data_9;
    assign token_9_7 = token_out_vec_9[6];
    assign dep_chan_vld_9_11 = out_chan_dep_vld_vec_9[7];
    assign dep_chan_data_9_11 = out_chan_dep_data_9;
    assign token_9_11 = token_out_vec_9[7];
    assign dep_chan_vld_9_12 = out_chan_dep_vld_vec_9[8];
    assign dep_chan_data_9_12 = out_chan_dep_data_9;
    assign token_9_12 = token_out_vec_9[8];
    assign dep_chan_vld_9_13 = out_chan_dep_vld_vec_9[9];
    assign dep_chan_data_9_13 = out_chan_dep_data_9;
    assign token_9_13 = token_out_vec_9[9];
    assign dep_chan_vld_9_14 = out_chan_dep_vld_vec_9[10];
    assign dep_chan_data_9_14 = out_chan_dep_data_9;
    assign token_9_14 = token_out_vec_9[10];
    assign dep_chan_vld_9_15 = out_chan_dep_vld_vec_9[11];
    assign dep_chan_data_9_15 = out_chan_dep_data_9;
    assign token_9_15 = token_out_vec_9[11];
    assign dep_chan_vld_9_16 = out_chan_dep_vld_vec_9[12];
    assign dep_chan_data_9_16 = out_chan_dep_data_9;
    assign token_9_16 = token_out_vec_9[12];
    assign dep_chan_vld_9_17 = out_chan_dep_vld_vec_9[13];
    assign dep_chan_data_9_17 = out_chan_dep_data_9;
    assign token_9_17 = token_out_vec_9[13];
    assign dep_chan_vld_9_18 = out_chan_dep_vld_vec_9[14];
    assign dep_chan_data_9_18 = out_chan_dep_data_9;
    assign token_9_18 = token_out_vec_9[14];
    assign dep_chan_vld_9_19 = out_chan_dep_vld_vec_9[15];
    assign dep_chan_data_9_19 = out_chan_dep_data_9;
    assign token_9_19 = token_out_vec_9[15];
    assign dep_chan_vld_9_20 = out_chan_dep_vld_vec_9[16];
    assign dep_chan_data_9_20 = out_chan_dep_data_9;
    assign token_9_20 = token_out_vec_9[16];
    assign dep_chan_vld_9_21 = out_chan_dep_vld_vec_9[17];
    assign dep_chan_data_9_21 = out_chan_dep_data_9;
    assign token_9_21 = token_out_vec_9[17];
    assign dep_chan_vld_9_22 = out_chan_dep_vld_vec_9[18];
    assign dep_chan_data_9_22 = out_chan_dep_data_9;
    assign token_9_22 = token_out_vec_9[18];
    assign dep_chan_vld_9_23 = out_chan_dep_vld_vec_9[19];
    assign dep_chan_data_9_23 = out_chan_dep_data_9;
    assign token_9_23 = token_out_vec_9[19];
    assign dep_chan_vld_9_24 = out_chan_dep_vld_vec_9[20];
    assign dep_chan_data_9_24 = out_chan_dep_data_9;
    assign token_9_24 = token_out_vec_9[20];
    assign dep_chan_vld_9_25 = out_chan_dep_vld_vec_9[21];
    assign dep_chan_data_9_25 = out_chan_dep_data_9;
    assign token_9_25 = token_out_vec_9[21];
    assign dep_chan_vld_9_26 = out_chan_dep_vld_vec_9[22];
    assign dep_chan_data_9_26 = out_chan_dep_data_9;
    assign token_9_26 = token_out_vec_9[22];
    assign dep_chan_vld_9_27 = out_chan_dep_vld_vec_9[23];
    assign dep_chan_data_9_27 = out_chan_dep_data_9;
    assign token_9_27 = token_out_vec_9[23];
    assign dep_chan_vld_9_28 = out_chan_dep_vld_vec_9[24];
    assign dep_chan_data_9_28 = out_chan_dep_data_9;
    assign token_9_28 = token_out_vec_9[24];
    assign dep_chan_vld_9_29 = out_chan_dep_vld_vec_9[25];
    assign dep_chan_data_9_29 = out_chan_dep_data_9;
    assign token_9_29 = token_out_vec_9[25];
    assign dep_chan_vld_9_30 = out_chan_dep_vld_vec_9[26];
    assign dep_chan_data_9_30 = out_chan_dep_data_9;
    assign token_9_30 = token_out_vec_9[26];
    assign dep_chan_vld_9_31 = out_chan_dep_vld_vec_9[27];
    assign dep_chan_data_9_31 = out_chan_dep_data_9;
    assign token_9_31 = token_out_vec_9[27];
    assign dep_chan_vld_9_32 = out_chan_dep_vld_vec_9[28];
    assign dep_chan_data_9_32 = out_chan_dep_data_9;
    assign token_9_32 = token_out_vec_9[28];
    assign dep_chan_vld_9_33 = out_chan_dep_vld_vec_9[29];
    assign dep_chan_data_9_33 = out_chan_dep_data_9;
    assign token_9_33 = token_out_vec_9[29];
    assign dep_chan_vld_9_34 = out_chan_dep_vld_vec_9[30];
    assign dep_chan_data_9_34 = out_chan_dep_data_9;
    assign token_9_34 = token_out_vec_9[30];
    assign dep_chan_vld_9_35 = out_chan_dep_vld_vec_9[31];
    assign dep_chan_data_9_35 = out_chan_dep_data_9;
    assign token_9_35 = token_out_vec_9[31];
    assign dep_chan_vld_9_36 = out_chan_dep_vld_vec_9[32];
    assign dep_chan_data_9_36 = out_chan_dep_data_9;
    assign token_9_36 = token_out_vec_9[32];

    // Process: ProcessingElement_5_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 10, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_10 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_10),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_10),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_10),
        .token_in_vec(token_in_vec_10),
        .dl_detect_in(dl_detect_out),
        .origin(origin[10]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_10),
        .out_chan_dep_data(out_chan_dep_data_10),
        .token_out_vec(token_out_vec_10),
        .dl_detect_out(dl_in_vec[10]));

    assign proc_10_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_4_blk_n) | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_4_blk_n) | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_WriteC_Flattened_fu_179.cPipes_4_blk_n);
    assign proc_10_data_PIPO_blk[0] = 1'b0;
    assign proc_10_start_FIFO_blk[0] = 1'b0;
    assign proc_10_TLF_FIFO_blk[0] = 1'b0;
    assign proc_10_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_10_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_10[0] = dl_detect_out ? proc_dep_vld_vec_10_reg[0] : (proc_10_data_FIFO_blk[0] | proc_10_data_PIPO_blk[0] | proc_10_start_FIFO_blk[0] | proc_10_TLF_FIFO_blk[0] | proc_10_input_sync_blk[0] | proc_10_output_sync_blk[0]);
    assign proc_10_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_5_blk_n) | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_5_blk_n) | (~ProcessingElement_5_U0.grp_ProcessingElement_5_Pipeline_WriteC_Flattened_fu_179.cPipes_5_blk_n);
    assign proc_10_data_PIPO_blk[1] = 1'b0;
    assign proc_10_start_FIFO_blk[1] = 1'b0;
    assign proc_10_TLF_FIFO_blk[1] = 1'b0;
    assign proc_10_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_10_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_10[1] = dl_detect_out ? proc_dep_vld_vec_10_reg[1] : (proc_10_data_FIFO_blk[1] | proc_10_data_PIPO_blk[1] | proc_10_start_FIFO_blk[1] | proc_10_TLF_FIFO_blk[1] | proc_10_input_sync_blk[1] | proc_10_output_sync_blk[1]);
    assign proc_10_data_FIFO_blk[2] = 1'b0;
    assign proc_10_data_PIPO_blk[2] = 1'b0;
    assign proc_10_start_FIFO_blk[2] = 1'b0;
    assign proc_10_TLF_FIFO_blk[2] = 1'b0;
    assign proc_10_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_10_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_10[2] = dl_detect_out ? proc_dep_vld_vec_10_reg[2] : (proc_10_data_FIFO_blk[2] | proc_10_data_PIPO_blk[2] | proc_10_start_FIFO_blk[2] | proc_10_TLF_FIFO_blk[2] | proc_10_input_sync_blk[2] | proc_10_output_sync_blk[2]);
    assign proc_10_data_FIFO_blk[3] = 1'b0;
    assign proc_10_data_PIPO_blk[3] = 1'b0;
    assign proc_10_start_FIFO_blk[3] = 1'b0;
    assign proc_10_TLF_FIFO_blk[3] = 1'b0;
    assign proc_10_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_10_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_10[3] = dl_detect_out ? proc_dep_vld_vec_10_reg[3] : (proc_10_data_FIFO_blk[3] | proc_10_data_PIPO_blk[3] | proc_10_start_FIFO_blk[3] | proc_10_TLF_FIFO_blk[3] | proc_10_input_sync_blk[3] | proc_10_output_sync_blk[3]);
    assign proc_10_data_FIFO_blk[4] = 1'b0;
    assign proc_10_data_PIPO_blk[4] = 1'b0;
    assign proc_10_start_FIFO_blk[4] = 1'b0;
    assign proc_10_TLF_FIFO_blk[4] = 1'b0;
    assign proc_10_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_10_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_10[4] = dl_detect_out ? proc_dep_vld_vec_10_reg[4] : (proc_10_data_FIFO_blk[4] | proc_10_data_PIPO_blk[4] | proc_10_start_FIFO_blk[4] | proc_10_TLF_FIFO_blk[4] | proc_10_input_sync_blk[4] | proc_10_output_sync_blk[4]);
    assign proc_10_data_FIFO_blk[5] = 1'b0;
    assign proc_10_data_PIPO_blk[5] = 1'b0;
    assign proc_10_start_FIFO_blk[5] = 1'b0;
    assign proc_10_TLF_FIFO_blk[5] = 1'b0;
    assign proc_10_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_10_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_10[5] = dl_detect_out ? proc_dep_vld_vec_10_reg[5] : (proc_10_data_FIFO_blk[5] | proc_10_data_PIPO_blk[5] | proc_10_start_FIFO_blk[5] | proc_10_TLF_FIFO_blk[5] | proc_10_input_sync_blk[5] | proc_10_output_sync_blk[5]);
    assign proc_10_data_FIFO_blk[6] = 1'b0;
    assign proc_10_data_PIPO_blk[6] = 1'b0;
    assign proc_10_start_FIFO_blk[6] = 1'b0;
    assign proc_10_TLF_FIFO_blk[6] = 1'b0;
    assign proc_10_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_10_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_10[6] = dl_detect_out ? proc_dep_vld_vec_10_reg[6] : (proc_10_data_FIFO_blk[6] | proc_10_data_PIPO_blk[6] | proc_10_start_FIFO_blk[6] | proc_10_TLF_FIFO_blk[6] | proc_10_input_sync_blk[6] | proc_10_output_sync_blk[6]);
    assign proc_10_data_FIFO_blk[7] = 1'b0;
    assign proc_10_data_PIPO_blk[7] = 1'b0;
    assign proc_10_start_FIFO_blk[7] = 1'b0;
    assign proc_10_TLF_FIFO_blk[7] = 1'b0;
    assign proc_10_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_10_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_10[7] = dl_detect_out ? proc_dep_vld_vec_10_reg[7] : (proc_10_data_FIFO_blk[7] | proc_10_data_PIPO_blk[7] | proc_10_start_FIFO_blk[7] | proc_10_TLF_FIFO_blk[7] | proc_10_input_sync_blk[7] | proc_10_output_sync_blk[7]);
    assign proc_10_data_FIFO_blk[8] = 1'b0;
    assign proc_10_data_PIPO_blk[8] = 1'b0;
    assign proc_10_start_FIFO_blk[8] = 1'b0;
    assign proc_10_TLF_FIFO_blk[8] = 1'b0;
    assign proc_10_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_10_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_10[8] = dl_detect_out ? proc_dep_vld_vec_10_reg[8] : (proc_10_data_FIFO_blk[8] | proc_10_data_PIPO_blk[8] | proc_10_start_FIFO_blk[8] | proc_10_TLF_FIFO_blk[8] | proc_10_input_sync_blk[8] | proc_10_output_sync_blk[8]);
    assign proc_10_data_FIFO_blk[9] = 1'b0;
    assign proc_10_data_PIPO_blk[9] = 1'b0;
    assign proc_10_start_FIFO_blk[9] = 1'b0;
    assign proc_10_TLF_FIFO_blk[9] = 1'b0;
    assign proc_10_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_10_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_10[9] = dl_detect_out ? proc_dep_vld_vec_10_reg[9] : (proc_10_data_FIFO_blk[9] | proc_10_data_PIPO_blk[9] | proc_10_start_FIFO_blk[9] | proc_10_TLF_FIFO_blk[9] | proc_10_input_sync_blk[9] | proc_10_output_sync_blk[9]);
    assign proc_10_data_FIFO_blk[10] = 1'b0;
    assign proc_10_data_PIPO_blk[10] = 1'b0;
    assign proc_10_start_FIFO_blk[10] = 1'b0;
    assign proc_10_TLF_FIFO_blk[10] = 1'b0;
    assign proc_10_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_10_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_10[10] = dl_detect_out ? proc_dep_vld_vec_10_reg[10] : (proc_10_data_FIFO_blk[10] | proc_10_data_PIPO_blk[10] | proc_10_start_FIFO_blk[10] | proc_10_TLF_FIFO_blk[10] | proc_10_input_sync_blk[10] | proc_10_output_sync_blk[10]);
    assign proc_10_data_FIFO_blk[11] = 1'b0;
    assign proc_10_data_PIPO_blk[11] = 1'b0;
    assign proc_10_start_FIFO_blk[11] = 1'b0;
    assign proc_10_TLF_FIFO_blk[11] = 1'b0;
    assign proc_10_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_10_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_10[11] = dl_detect_out ? proc_dep_vld_vec_10_reg[11] : (proc_10_data_FIFO_blk[11] | proc_10_data_PIPO_blk[11] | proc_10_start_FIFO_blk[11] | proc_10_TLF_FIFO_blk[11] | proc_10_input_sync_blk[11] | proc_10_output_sync_blk[11]);
    assign proc_10_data_FIFO_blk[12] = 1'b0;
    assign proc_10_data_PIPO_blk[12] = 1'b0;
    assign proc_10_start_FIFO_blk[12] = 1'b0;
    assign proc_10_TLF_FIFO_blk[12] = 1'b0;
    assign proc_10_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_10_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_10[12] = dl_detect_out ? proc_dep_vld_vec_10_reg[12] : (proc_10_data_FIFO_blk[12] | proc_10_data_PIPO_blk[12] | proc_10_start_FIFO_blk[12] | proc_10_TLF_FIFO_blk[12] | proc_10_input_sync_blk[12] | proc_10_output_sync_blk[12]);
    assign proc_10_data_FIFO_blk[13] = 1'b0;
    assign proc_10_data_PIPO_blk[13] = 1'b0;
    assign proc_10_start_FIFO_blk[13] = 1'b0;
    assign proc_10_TLF_FIFO_blk[13] = 1'b0;
    assign proc_10_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_10_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_10[13] = dl_detect_out ? proc_dep_vld_vec_10_reg[13] : (proc_10_data_FIFO_blk[13] | proc_10_data_PIPO_blk[13] | proc_10_start_FIFO_blk[13] | proc_10_TLF_FIFO_blk[13] | proc_10_input_sync_blk[13] | proc_10_output_sync_blk[13]);
    assign proc_10_data_FIFO_blk[14] = 1'b0;
    assign proc_10_data_PIPO_blk[14] = 1'b0;
    assign proc_10_start_FIFO_blk[14] = 1'b0;
    assign proc_10_TLF_FIFO_blk[14] = 1'b0;
    assign proc_10_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_10_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_10[14] = dl_detect_out ? proc_dep_vld_vec_10_reg[14] : (proc_10_data_FIFO_blk[14] | proc_10_data_PIPO_blk[14] | proc_10_start_FIFO_blk[14] | proc_10_TLF_FIFO_blk[14] | proc_10_input_sync_blk[14] | proc_10_output_sync_blk[14]);
    assign proc_10_data_FIFO_blk[15] = 1'b0;
    assign proc_10_data_PIPO_blk[15] = 1'b0;
    assign proc_10_start_FIFO_blk[15] = 1'b0;
    assign proc_10_TLF_FIFO_blk[15] = 1'b0;
    assign proc_10_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_10_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_10[15] = dl_detect_out ? proc_dep_vld_vec_10_reg[15] : (proc_10_data_FIFO_blk[15] | proc_10_data_PIPO_blk[15] | proc_10_start_FIFO_blk[15] | proc_10_TLF_FIFO_blk[15] | proc_10_input_sync_blk[15] | proc_10_output_sync_blk[15]);
    assign proc_10_data_FIFO_blk[16] = 1'b0;
    assign proc_10_data_PIPO_blk[16] = 1'b0;
    assign proc_10_start_FIFO_blk[16] = 1'b0;
    assign proc_10_TLF_FIFO_blk[16] = 1'b0;
    assign proc_10_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_10_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_10[16] = dl_detect_out ? proc_dep_vld_vec_10_reg[16] : (proc_10_data_FIFO_blk[16] | proc_10_data_PIPO_blk[16] | proc_10_start_FIFO_blk[16] | proc_10_TLF_FIFO_blk[16] | proc_10_input_sync_blk[16] | proc_10_output_sync_blk[16]);
    assign proc_10_data_FIFO_blk[17] = 1'b0;
    assign proc_10_data_PIPO_blk[17] = 1'b0;
    assign proc_10_start_FIFO_blk[17] = 1'b0;
    assign proc_10_TLF_FIFO_blk[17] = 1'b0;
    assign proc_10_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_10_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_10[17] = dl_detect_out ? proc_dep_vld_vec_10_reg[17] : (proc_10_data_FIFO_blk[17] | proc_10_data_PIPO_blk[17] | proc_10_start_FIFO_blk[17] | proc_10_TLF_FIFO_blk[17] | proc_10_input_sync_blk[17] | proc_10_output_sync_blk[17]);
    assign proc_10_data_FIFO_blk[18] = 1'b0;
    assign proc_10_data_PIPO_blk[18] = 1'b0;
    assign proc_10_start_FIFO_blk[18] = 1'b0;
    assign proc_10_TLF_FIFO_blk[18] = 1'b0;
    assign proc_10_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_10_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_10[18] = dl_detect_out ? proc_dep_vld_vec_10_reg[18] : (proc_10_data_FIFO_blk[18] | proc_10_data_PIPO_blk[18] | proc_10_start_FIFO_blk[18] | proc_10_TLF_FIFO_blk[18] | proc_10_input_sync_blk[18] | proc_10_output_sync_blk[18]);
    assign proc_10_data_FIFO_blk[19] = 1'b0;
    assign proc_10_data_PIPO_blk[19] = 1'b0;
    assign proc_10_start_FIFO_blk[19] = 1'b0;
    assign proc_10_TLF_FIFO_blk[19] = 1'b0;
    assign proc_10_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_10_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_10[19] = dl_detect_out ? proc_dep_vld_vec_10_reg[19] : (proc_10_data_FIFO_blk[19] | proc_10_data_PIPO_blk[19] | proc_10_start_FIFO_blk[19] | proc_10_TLF_FIFO_blk[19] | proc_10_input_sync_blk[19] | proc_10_output_sync_blk[19]);
    assign proc_10_data_FIFO_blk[20] = 1'b0;
    assign proc_10_data_PIPO_blk[20] = 1'b0;
    assign proc_10_start_FIFO_blk[20] = 1'b0;
    assign proc_10_TLF_FIFO_blk[20] = 1'b0;
    assign proc_10_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_10_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_10[20] = dl_detect_out ? proc_dep_vld_vec_10_reg[20] : (proc_10_data_FIFO_blk[20] | proc_10_data_PIPO_blk[20] | proc_10_start_FIFO_blk[20] | proc_10_TLF_FIFO_blk[20] | proc_10_input_sync_blk[20] | proc_10_output_sync_blk[20]);
    assign proc_10_data_FIFO_blk[21] = 1'b0;
    assign proc_10_data_PIPO_blk[21] = 1'b0;
    assign proc_10_start_FIFO_blk[21] = 1'b0;
    assign proc_10_TLF_FIFO_blk[21] = 1'b0;
    assign proc_10_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_10_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_10[21] = dl_detect_out ? proc_dep_vld_vec_10_reg[21] : (proc_10_data_FIFO_blk[21] | proc_10_data_PIPO_blk[21] | proc_10_start_FIFO_blk[21] | proc_10_TLF_FIFO_blk[21] | proc_10_input_sync_blk[21] | proc_10_output_sync_blk[21]);
    assign proc_10_data_FIFO_blk[22] = 1'b0;
    assign proc_10_data_PIPO_blk[22] = 1'b0;
    assign proc_10_start_FIFO_blk[22] = 1'b0;
    assign proc_10_TLF_FIFO_blk[22] = 1'b0;
    assign proc_10_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_10_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_10[22] = dl_detect_out ? proc_dep_vld_vec_10_reg[22] : (proc_10_data_FIFO_blk[22] | proc_10_data_PIPO_blk[22] | proc_10_start_FIFO_blk[22] | proc_10_TLF_FIFO_blk[22] | proc_10_input_sync_blk[22] | proc_10_output_sync_blk[22]);
    assign proc_10_data_FIFO_blk[23] = 1'b0;
    assign proc_10_data_PIPO_blk[23] = 1'b0;
    assign proc_10_start_FIFO_blk[23] = 1'b0;
    assign proc_10_TLF_FIFO_blk[23] = 1'b0;
    assign proc_10_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_10_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_10[23] = dl_detect_out ? proc_dep_vld_vec_10_reg[23] : (proc_10_data_FIFO_blk[23] | proc_10_data_PIPO_blk[23] | proc_10_start_FIFO_blk[23] | proc_10_TLF_FIFO_blk[23] | proc_10_input_sync_blk[23] | proc_10_output_sync_blk[23]);
    assign proc_10_data_FIFO_blk[24] = 1'b0;
    assign proc_10_data_PIPO_blk[24] = 1'b0;
    assign proc_10_start_FIFO_blk[24] = 1'b0;
    assign proc_10_TLF_FIFO_blk[24] = 1'b0;
    assign proc_10_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_10_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_10[24] = dl_detect_out ? proc_dep_vld_vec_10_reg[24] : (proc_10_data_FIFO_blk[24] | proc_10_data_PIPO_blk[24] | proc_10_start_FIFO_blk[24] | proc_10_TLF_FIFO_blk[24] | proc_10_input_sync_blk[24] | proc_10_output_sync_blk[24]);
    assign proc_10_data_FIFO_blk[25] = 1'b0;
    assign proc_10_data_PIPO_blk[25] = 1'b0;
    assign proc_10_start_FIFO_blk[25] = 1'b0;
    assign proc_10_TLF_FIFO_blk[25] = 1'b0;
    assign proc_10_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_10_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_10[25] = dl_detect_out ? proc_dep_vld_vec_10_reg[25] : (proc_10_data_FIFO_blk[25] | proc_10_data_PIPO_blk[25] | proc_10_start_FIFO_blk[25] | proc_10_TLF_FIFO_blk[25] | proc_10_input_sync_blk[25] | proc_10_output_sync_blk[25]);
    assign proc_10_data_FIFO_blk[26] = 1'b0;
    assign proc_10_data_PIPO_blk[26] = 1'b0;
    assign proc_10_start_FIFO_blk[26] = 1'b0;
    assign proc_10_TLF_FIFO_blk[26] = 1'b0;
    assign proc_10_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_10_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_10[26] = dl_detect_out ? proc_dep_vld_vec_10_reg[26] : (proc_10_data_FIFO_blk[26] | proc_10_data_PIPO_blk[26] | proc_10_start_FIFO_blk[26] | proc_10_TLF_FIFO_blk[26] | proc_10_input_sync_blk[26] | proc_10_output_sync_blk[26]);
    assign proc_10_data_FIFO_blk[27] = 1'b0;
    assign proc_10_data_PIPO_blk[27] = 1'b0;
    assign proc_10_start_FIFO_blk[27] = 1'b0;
    assign proc_10_TLF_FIFO_blk[27] = 1'b0;
    assign proc_10_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_10_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_10[27] = dl_detect_out ? proc_dep_vld_vec_10_reg[27] : (proc_10_data_FIFO_blk[27] | proc_10_data_PIPO_blk[27] | proc_10_start_FIFO_blk[27] | proc_10_TLF_FIFO_blk[27] | proc_10_input_sync_blk[27] | proc_10_output_sync_blk[27]);
    assign proc_10_data_FIFO_blk[28] = 1'b0;
    assign proc_10_data_PIPO_blk[28] = 1'b0;
    assign proc_10_start_FIFO_blk[28] = 1'b0;
    assign proc_10_TLF_FIFO_blk[28] = 1'b0;
    assign proc_10_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_10_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_10[28] = dl_detect_out ? proc_dep_vld_vec_10_reg[28] : (proc_10_data_FIFO_blk[28] | proc_10_data_PIPO_blk[28] | proc_10_start_FIFO_blk[28] | proc_10_TLF_FIFO_blk[28] | proc_10_input_sync_blk[28] | proc_10_output_sync_blk[28]);
    assign proc_10_data_FIFO_blk[29] = 1'b0;
    assign proc_10_data_PIPO_blk[29] = 1'b0;
    assign proc_10_start_FIFO_blk[29] = 1'b0;
    assign proc_10_TLF_FIFO_blk[29] = 1'b0;
    assign proc_10_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_10_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_10[29] = dl_detect_out ? proc_dep_vld_vec_10_reg[29] : (proc_10_data_FIFO_blk[29] | proc_10_data_PIPO_blk[29] | proc_10_start_FIFO_blk[29] | proc_10_TLF_FIFO_blk[29] | proc_10_input_sync_blk[29] | proc_10_output_sync_blk[29]);
    assign proc_10_data_FIFO_blk[30] = 1'b0;
    assign proc_10_data_PIPO_blk[30] = 1'b0;
    assign proc_10_start_FIFO_blk[30] = 1'b0;
    assign proc_10_TLF_FIFO_blk[30] = 1'b0;
    assign proc_10_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_10_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_10[30] = dl_detect_out ? proc_dep_vld_vec_10_reg[30] : (proc_10_data_FIFO_blk[30] | proc_10_data_PIPO_blk[30] | proc_10_start_FIFO_blk[30] | proc_10_TLF_FIFO_blk[30] | proc_10_input_sync_blk[30] | proc_10_output_sync_blk[30]);
    assign proc_10_data_FIFO_blk[31] = 1'b0;
    assign proc_10_data_PIPO_blk[31] = 1'b0;
    assign proc_10_start_FIFO_blk[31] = 1'b0;
    assign proc_10_TLF_FIFO_blk[31] = 1'b0;
    assign proc_10_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_10_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_10[31] = dl_detect_out ? proc_dep_vld_vec_10_reg[31] : (proc_10_data_FIFO_blk[31] | proc_10_data_PIPO_blk[31] | proc_10_start_FIFO_blk[31] | proc_10_TLF_FIFO_blk[31] | proc_10_input_sync_blk[31] | proc_10_output_sync_blk[31]);
    assign proc_10_data_FIFO_blk[32] = 1'b0;
    assign proc_10_data_PIPO_blk[32] = 1'b0;
    assign proc_10_start_FIFO_blk[32] = 1'b0;
    assign proc_10_TLF_FIFO_blk[32] = 1'b0;
    assign proc_10_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_5_U0_ap_ready & ProcessingElement_5_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_10_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_10[32] = dl_detect_out ? proc_dep_vld_vec_10_reg[32] : (proc_10_data_FIFO_blk[32] | proc_10_data_PIPO_blk[32] | proc_10_start_FIFO_blk[32] | proc_10_TLF_FIFO_blk[32] | proc_10_input_sync_blk[32] | proc_10_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_10_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_10_reg <= proc_dep_vld_vec_10;
        end
    end
    assign in_chan_dep_vld_vec_10[0] = dep_chan_vld_0_10;
    assign in_chan_dep_data_vec_10[39 : 0] = dep_chan_data_0_10;
    assign token_in_vec_10[0] = token_0_10;
    assign in_chan_dep_vld_vec_10[1] = dep_chan_vld_1_10;
    assign in_chan_dep_data_vec_10[79 : 40] = dep_chan_data_1_10;
    assign token_in_vec_10[1] = token_1_10;
    assign in_chan_dep_vld_vec_10[2] = dep_chan_vld_3_10;
    assign in_chan_dep_data_vec_10[119 : 80] = dep_chan_data_3_10;
    assign token_in_vec_10[2] = token_3_10;
    assign in_chan_dep_vld_vec_10[3] = dep_chan_vld_6_10;
    assign in_chan_dep_data_vec_10[159 : 120] = dep_chan_data_6_10;
    assign token_in_vec_10[3] = token_6_10;
    assign in_chan_dep_vld_vec_10[4] = dep_chan_vld_7_10;
    assign in_chan_dep_data_vec_10[199 : 160] = dep_chan_data_7_10;
    assign token_in_vec_10[4] = token_7_10;
    assign in_chan_dep_vld_vec_10[5] = dep_chan_vld_8_10;
    assign in_chan_dep_data_vec_10[239 : 200] = dep_chan_data_8_10;
    assign token_in_vec_10[5] = token_8_10;
    assign in_chan_dep_vld_vec_10[6] = dep_chan_vld_9_10;
    assign in_chan_dep_data_vec_10[279 : 240] = dep_chan_data_9_10;
    assign token_in_vec_10[6] = token_9_10;
    assign in_chan_dep_vld_vec_10[7] = dep_chan_vld_11_10;
    assign in_chan_dep_data_vec_10[319 : 280] = dep_chan_data_11_10;
    assign token_in_vec_10[7] = token_11_10;
    assign in_chan_dep_vld_vec_10[8] = dep_chan_vld_12_10;
    assign in_chan_dep_data_vec_10[359 : 320] = dep_chan_data_12_10;
    assign token_in_vec_10[8] = token_12_10;
    assign in_chan_dep_vld_vec_10[9] = dep_chan_vld_13_10;
    assign in_chan_dep_data_vec_10[399 : 360] = dep_chan_data_13_10;
    assign token_in_vec_10[9] = token_13_10;
    assign in_chan_dep_vld_vec_10[10] = dep_chan_vld_14_10;
    assign in_chan_dep_data_vec_10[439 : 400] = dep_chan_data_14_10;
    assign token_in_vec_10[10] = token_14_10;
    assign in_chan_dep_vld_vec_10[11] = dep_chan_vld_15_10;
    assign in_chan_dep_data_vec_10[479 : 440] = dep_chan_data_15_10;
    assign token_in_vec_10[11] = token_15_10;
    assign in_chan_dep_vld_vec_10[12] = dep_chan_vld_16_10;
    assign in_chan_dep_data_vec_10[519 : 480] = dep_chan_data_16_10;
    assign token_in_vec_10[12] = token_16_10;
    assign in_chan_dep_vld_vec_10[13] = dep_chan_vld_17_10;
    assign in_chan_dep_data_vec_10[559 : 520] = dep_chan_data_17_10;
    assign token_in_vec_10[13] = token_17_10;
    assign in_chan_dep_vld_vec_10[14] = dep_chan_vld_18_10;
    assign in_chan_dep_data_vec_10[599 : 560] = dep_chan_data_18_10;
    assign token_in_vec_10[14] = token_18_10;
    assign in_chan_dep_vld_vec_10[15] = dep_chan_vld_19_10;
    assign in_chan_dep_data_vec_10[639 : 600] = dep_chan_data_19_10;
    assign token_in_vec_10[15] = token_19_10;
    assign in_chan_dep_vld_vec_10[16] = dep_chan_vld_20_10;
    assign in_chan_dep_data_vec_10[679 : 640] = dep_chan_data_20_10;
    assign token_in_vec_10[16] = token_20_10;
    assign in_chan_dep_vld_vec_10[17] = dep_chan_vld_21_10;
    assign in_chan_dep_data_vec_10[719 : 680] = dep_chan_data_21_10;
    assign token_in_vec_10[17] = token_21_10;
    assign in_chan_dep_vld_vec_10[18] = dep_chan_vld_22_10;
    assign in_chan_dep_data_vec_10[759 : 720] = dep_chan_data_22_10;
    assign token_in_vec_10[18] = token_22_10;
    assign in_chan_dep_vld_vec_10[19] = dep_chan_vld_23_10;
    assign in_chan_dep_data_vec_10[799 : 760] = dep_chan_data_23_10;
    assign token_in_vec_10[19] = token_23_10;
    assign in_chan_dep_vld_vec_10[20] = dep_chan_vld_24_10;
    assign in_chan_dep_data_vec_10[839 : 800] = dep_chan_data_24_10;
    assign token_in_vec_10[20] = token_24_10;
    assign in_chan_dep_vld_vec_10[21] = dep_chan_vld_25_10;
    assign in_chan_dep_data_vec_10[879 : 840] = dep_chan_data_25_10;
    assign token_in_vec_10[21] = token_25_10;
    assign in_chan_dep_vld_vec_10[22] = dep_chan_vld_26_10;
    assign in_chan_dep_data_vec_10[919 : 880] = dep_chan_data_26_10;
    assign token_in_vec_10[22] = token_26_10;
    assign in_chan_dep_vld_vec_10[23] = dep_chan_vld_27_10;
    assign in_chan_dep_data_vec_10[959 : 920] = dep_chan_data_27_10;
    assign token_in_vec_10[23] = token_27_10;
    assign in_chan_dep_vld_vec_10[24] = dep_chan_vld_28_10;
    assign in_chan_dep_data_vec_10[999 : 960] = dep_chan_data_28_10;
    assign token_in_vec_10[24] = token_28_10;
    assign in_chan_dep_vld_vec_10[25] = dep_chan_vld_29_10;
    assign in_chan_dep_data_vec_10[1039 : 1000] = dep_chan_data_29_10;
    assign token_in_vec_10[25] = token_29_10;
    assign in_chan_dep_vld_vec_10[26] = dep_chan_vld_30_10;
    assign in_chan_dep_data_vec_10[1079 : 1040] = dep_chan_data_30_10;
    assign token_in_vec_10[26] = token_30_10;
    assign in_chan_dep_vld_vec_10[27] = dep_chan_vld_31_10;
    assign in_chan_dep_data_vec_10[1119 : 1080] = dep_chan_data_31_10;
    assign token_in_vec_10[27] = token_31_10;
    assign in_chan_dep_vld_vec_10[28] = dep_chan_vld_32_10;
    assign in_chan_dep_data_vec_10[1159 : 1120] = dep_chan_data_32_10;
    assign token_in_vec_10[28] = token_32_10;
    assign in_chan_dep_vld_vec_10[29] = dep_chan_vld_33_10;
    assign in_chan_dep_data_vec_10[1199 : 1160] = dep_chan_data_33_10;
    assign token_in_vec_10[29] = token_33_10;
    assign in_chan_dep_vld_vec_10[30] = dep_chan_vld_34_10;
    assign in_chan_dep_data_vec_10[1239 : 1200] = dep_chan_data_34_10;
    assign token_in_vec_10[30] = token_34_10;
    assign in_chan_dep_vld_vec_10[31] = dep_chan_vld_35_10;
    assign in_chan_dep_data_vec_10[1279 : 1240] = dep_chan_data_35_10;
    assign token_in_vec_10[31] = token_35_10;
    assign in_chan_dep_vld_vec_10[32] = dep_chan_vld_36_10;
    assign in_chan_dep_data_vec_10[1319 : 1280] = dep_chan_data_36_10;
    assign token_in_vec_10[32] = token_36_10;
    assign dep_chan_vld_10_9 = out_chan_dep_vld_vec_10[0];
    assign dep_chan_data_10_9 = out_chan_dep_data_10;
    assign token_10_9 = token_out_vec_10[0];
    assign dep_chan_vld_10_11 = out_chan_dep_vld_vec_10[1];
    assign dep_chan_data_10_11 = out_chan_dep_data_10;
    assign token_10_11 = token_out_vec_10[1];
    assign dep_chan_vld_10_0 = out_chan_dep_vld_vec_10[2];
    assign dep_chan_data_10_0 = out_chan_dep_data_10;
    assign token_10_0 = token_out_vec_10[2];
    assign dep_chan_vld_10_1 = out_chan_dep_vld_vec_10[3];
    assign dep_chan_data_10_1 = out_chan_dep_data_10;
    assign token_10_1 = token_out_vec_10[3];
    assign dep_chan_vld_10_3 = out_chan_dep_vld_vec_10[4];
    assign dep_chan_data_10_3 = out_chan_dep_data_10;
    assign token_10_3 = token_out_vec_10[4];
    assign dep_chan_vld_10_6 = out_chan_dep_vld_vec_10[5];
    assign dep_chan_data_10_6 = out_chan_dep_data_10;
    assign token_10_6 = token_out_vec_10[5];
    assign dep_chan_vld_10_7 = out_chan_dep_vld_vec_10[6];
    assign dep_chan_data_10_7 = out_chan_dep_data_10;
    assign token_10_7 = token_out_vec_10[6];
    assign dep_chan_vld_10_8 = out_chan_dep_vld_vec_10[7];
    assign dep_chan_data_10_8 = out_chan_dep_data_10;
    assign token_10_8 = token_out_vec_10[7];
    assign dep_chan_vld_10_12 = out_chan_dep_vld_vec_10[8];
    assign dep_chan_data_10_12 = out_chan_dep_data_10;
    assign token_10_12 = token_out_vec_10[8];
    assign dep_chan_vld_10_13 = out_chan_dep_vld_vec_10[9];
    assign dep_chan_data_10_13 = out_chan_dep_data_10;
    assign token_10_13 = token_out_vec_10[9];
    assign dep_chan_vld_10_14 = out_chan_dep_vld_vec_10[10];
    assign dep_chan_data_10_14 = out_chan_dep_data_10;
    assign token_10_14 = token_out_vec_10[10];
    assign dep_chan_vld_10_15 = out_chan_dep_vld_vec_10[11];
    assign dep_chan_data_10_15 = out_chan_dep_data_10;
    assign token_10_15 = token_out_vec_10[11];
    assign dep_chan_vld_10_16 = out_chan_dep_vld_vec_10[12];
    assign dep_chan_data_10_16 = out_chan_dep_data_10;
    assign token_10_16 = token_out_vec_10[12];
    assign dep_chan_vld_10_17 = out_chan_dep_vld_vec_10[13];
    assign dep_chan_data_10_17 = out_chan_dep_data_10;
    assign token_10_17 = token_out_vec_10[13];
    assign dep_chan_vld_10_18 = out_chan_dep_vld_vec_10[14];
    assign dep_chan_data_10_18 = out_chan_dep_data_10;
    assign token_10_18 = token_out_vec_10[14];
    assign dep_chan_vld_10_19 = out_chan_dep_vld_vec_10[15];
    assign dep_chan_data_10_19 = out_chan_dep_data_10;
    assign token_10_19 = token_out_vec_10[15];
    assign dep_chan_vld_10_20 = out_chan_dep_vld_vec_10[16];
    assign dep_chan_data_10_20 = out_chan_dep_data_10;
    assign token_10_20 = token_out_vec_10[16];
    assign dep_chan_vld_10_21 = out_chan_dep_vld_vec_10[17];
    assign dep_chan_data_10_21 = out_chan_dep_data_10;
    assign token_10_21 = token_out_vec_10[17];
    assign dep_chan_vld_10_22 = out_chan_dep_vld_vec_10[18];
    assign dep_chan_data_10_22 = out_chan_dep_data_10;
    assign token_10_22 = token_out_vec_10[18];
    assign dep_chan_vld_10_23 = out_chan_dep_vld_vec_10[19];
    assign dep_chan_data_10_23 = out_chan_dep_data_10;
    assign token_10_23 = token_out_vec_10[19];
    assign dep_chan_vld_10_24 = out_chan_dep_vld_vec_10[20];
    assign dep_chan_data_10_24 = out_chan_dep_data_10;
    assign token_10_24 = token_out_vec_10[20];
    assign dep_chan_vld_10_25 = out_chan_dep_vld_vec_10[21];
    assign dep_chan_data_10_25 = out_chan_dep_data_10;
    assign token_10_25 = token_out_vec_10[21];
    assign dep_chan_vld_10_26 = out_chan_dep_vld_vec_10[22];
    assign dep_chan_data_10_26 = out_chan_dep_data_10;
    assign token_10_26 = token_out_vec_10[22];
    assign dep_chan_vld_10_27 = out_chan_dep_vld_vec_10[23];
    assign dep_chan_data_10_27 = out_chan_dep_data_10;
    assign token_10_27 = token_out_vec_10[23];
    assign dep_chan_vld_10_28 = out_chan_dep_vld_vec_10[24];
    assign dep_chan_data_10_28 = out_chan_dep_data_10;
    assign token_10_28 = token_out_vec_10[24];
    assign dep_chan_vld_10_29 = out_chan_dep_vld_vec_10[25];
    assign dep_chan_data_10_29 = out_chan_dep_data_10;
    assign token_10_29 = token_out_vec_10[25];
    assign dep_chan_vld_10_30 = out_chan_dep_vld_vec_10[26];
    assign dep_chan_data_10_30 = out_chan_dep_data_10;
    assign token_10_30 = token_out_vec_10[26];
    assign dep_chan_vld_10_31 = out_chan_dep_vld_vec_10[27];
    assign dep_chan_data_10_31 = out_chan_dep_data_10;
    assign token_10_31 = token_out_vec_10[27];
    assign dep_chan_vld_10_32 = out_chan_dep_vld_vec_10[28];
    assign dep_chan_data_10_32 = out_chan_dep_data_10;
    assign token_10_32 = token_out_vec_10[28];
    assign dep_chan_vld_10_33 = out_chan_dep_vld_vec_10[29];
    assign dep_chan_data_10_33 = out_chan_dep_data_10;
    assign token_10_33 = token_out_vec_10[29];
    assign dep_chan_vld_10_34 = out_chan_dep_vld_vec_10[30];
    assign dep_chan_data_10_34 = out_chan_dep_data_10;
    assign token_10_34 = token_out_vec_10[30];
    assign dep_chan_vld_10_35 = out_chan_dep_vld_vec_10[31];
    assign dep_chan_data_10_35 = out_chan_dep_data_10;
    assign token_10_35 = token_out_vec_10[31];
    assign dep_chan_vld_10_36 = out_chan_dep_vld_vec_10[32];
    assign dep_chan_data_10_36 = out_chan_dep_data_10;
    assign token_10_36 = token_out_vec_10[32];

    // Process: ProcessingElement_6_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 11, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_11 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_11),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_11),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_11),
        .token_in_vec(token_in_vec_11),
        .dl_detect_in(dl_detect_out),
        .origin(origin[11]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_11),
        .out_chan_dep_data(out_chan_dep_data_11),
        .token_out_vec(token_out_vec_11),
        .dl_detect_out(dl_in_vec[11]));

    assign proc_11_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_5_blk_n) | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_5_blk_n) | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_WriteC_Flattened_fu_179.cPipes_5_blk_n);
    assign proc_11_data_PIPO_blk[0] = 1'b0;
    assign proc_11_start_FIFO_blk[0] = 1'b0;
    assign proc_11_TLF_FIFO_blk[0] = 1'b0;
    assign proc_11_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_11_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_11[0] = dl_detect_out ? proc_dep_vld_vec_11_reg[0] : (proc_11_data_FIFO_blk[0] | proc_11_data_PIPO_blk[0] | proc_11_start_FIFO_blk[0] | proc_11_TLF_FIFO_blk[0] | proc_11_input_sync_blk[0] | proc_11_output_sync_blk[0]);
    assign proc_11_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_6_blk_n) | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_6_blk_n) | (~ProcessingElement_6_U0.grp_ProcessingElement_6_Pipeline_WriteC_Flattened_fu_179.cPipes_6_blk_n);
    assign proc_11_data_PIPO_blk[1] = 1'b0;
    assign proc_11_start_FIFO_blk[1] = 1'b0;
    assign proc_11_TLF_FIFO_blk[1] = 1'b0;
    assign proc_11_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_11_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_11[1] = dl_detect_out ? proc_dep_vld_vec_11_reg[1] : (proc_11_data_FIFO_blk[1] | proc_11_data_PIPO_blk[1] | proc_11_start_FIFO_blk[1] | proc_11_TLF_FIFO_blk[1] | proc_11_input_sync_blk[1] | proc_11_output_sync_blk[1]);
    assign proc_11_data_FIFO_blk[2] = 1'b0;
    assign proc_11_data_PIPO_blk[2] = 1'b0;
    assign proc_11_start_FIFO_blk[2] = 1'b0;
    assign proc_11_TLF_FIFO_blk[2] = 1'b0;
    assign proc_11_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_11_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_11[2] = dl_detect_out ? proc_dep_vld_vec_11_reg[2] : (proc_11_data_FIFO_blk[2] | proc_11_data_PIPO_blk[2] | proc_11_start_FIFO_blk[2] | proc_11_TLF_FIFO_blk[2] | proc_11_input_sync_blk[2] | proc_11_output_sync_blk[2]);
    assign proc_11_data_FIFO_blk[3] = 1'b0;
    assign proc_11_data_PIPO_blk[3] = 1'b0;
    assign proc_11_start_FIFO_blk[3] = 1'b0;
    assign proc_11_TLF_FIFO_blk[3] = 1'b0;
    assign proc_11_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_11_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_11[3] = dl_detect_out ? proc_dep_vld_vec_11_reg[3] : (proc_11_data_FIFO_blk[3] | proc_11_data_PIPO_blk[3] | proc_11_start_FIFO_blk[3] | proc_11_TLF_FIFO_blk[3] | proc_11_input_sync_blk[3] | proc_11_output_sync_blk[3]);
    assign proc_11_data_FIFO_blk[4] = 1'b0;
    assign proc_11_data_PIPO_blk[4] = 1'b0;
    assign proc_11_start_FIFO_blk[4] = 1'b0;
    assign proc_11_TLF_FIFO_blk[4] = 1'b0;
    assign proc_11_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_11_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_11[4] = dl_detect_out ? proc_dep_vld_vec_11_reg[4] : (proc_11_data_FIFO_blk[4] | proc_11_data_PIPO_blk[4] | proc_11_start_FIFO_blk[4] | proc_11_TLF_FIFO_blk[4] | proc_11_input_sync_blk[4] | proc_11_output_sync_blk[4]);
    assign proc_11_data_FIFO_blk[5] = 1'b0;
    assign proc_11_data_PIPO_blk[5] = 1'b0;
    assign proc_11_start_FIFO_blk[5] = 1'b0;
    assign proc_11_TLF_FIFO_blk[5] = 1'b0;
    assign proc_11_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_11_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_11[5] = dl_detect_out ? proc_dep_vld_vec_11_reg[5] : (proc_11_data_FIFO_blk[5] | proc_11_data_PIPO_blk[5] | proc_11_start_FIFO_blk[5] | proc_11_TLF_FIFO_blk[5] | proc_11_input_sync_blk[5] | proc_11_output_sync_blk[5]);
    assign proc_11_data_FIFO_blk[6] = 1'b0;
    assign proc_11_data_PIPO_blk[6] = 1'b0;
    assign proc_11_start_FIFO_blk[6] = 1'b0;
    assign proc_11_TLF_FIFO_blk[6] = 1'b0;
    assign proc_11_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_11_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_11[6] = dl_detect_out ? proc_dep_vld_vec_11_reg[6] : (proc_11_data_FIFO_blk[6] | proc_11_data_PIPO_blk[6] | proc_11_start_FIFO_blk[6] | proc_11_TLF_FIFO_blk[6] | proc_11_input_sync_blk[6] | proc_11_output_sync_blk[6]);
    assign proc_11_data_FIFO_blk[7] = 1'b0;
    assign proc_11_data_PIPO_blk[7] = 1'b0;
    assign proc_11_start_FIFO_blk[7] = 1'b0;
    assign proc_11_TLF_FIFO_blk[7] = 1'b0;
    assign proc_11_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_11_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_11[7] = dl_detect_out ? proc_dep_vld_vec_11_reg[7] : (proc_11_data_FIFO_blk[7] | proc_11_data_PIPO_blk[7] | proc_11_start_FIFO_blk[7] | proc_11_TLF_FIFO_blk[7] | proc_11_input_sync_blk[7] | proc_11_output_sync_blk[7]);
    assign proc_11_data_FIFO_blk[8] = 1'b0;
    assign proc_11_data_PIPO_blk[8] = 1'b0;
    assign proc_11_start_FIFO_blk[8] = 1'b0;
    assign proc_11_TLF_FIFO_blk[8] = 1'b0;
    assign proc_11_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_11_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_11[8] = dl_detect_out ? proc_dep_vld_vec_11_reg[8] : (proc_11_data_FIFO_blk[8] | proc_11_data_PIPO_blk[8] | proc_11_start_FIFO_blk[8] | proc_11_TLF_FIFO_blk[8] | proc_11_input_sync_blk[8] | proc_11_output_sync_blk[8]);
    assign proc_11_data_FIFO_blk[9] = 1'b0;
    assign proc_11_data_PIPO_blk[9] = 1'b0;
    assign proc_11_start_FIFO_blk[9] = 1'b0;
    assign proc_11_TLF_FIFO_blk[9] = 1'b0;
    assign proc_11_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_11_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_11[9] = dl_detect_out ? proc_dep_vld_vec_11_reg[9] : (proc_11_data_FIFO_blk[9] | proc_11_data_PIPO_blk[9] | proc_11_start_FIFO_blk[9] | proc_11_TLF_FIFO_blk[9] | proc_11_input_sync_blk[9] | proc_11_output_sync_blk[9]);
    assign proc_11_data_FIFO_blk[10] = 1'b0;
    assign proc_11_data_PIPO_blk[10] = 1'b0;
    assign proc_11_start_FIFO_blk[10] = 1'b0;
    assign proc_11_TLF_FIFO_blk[10] = 1'b0;
    assign proc_11_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_11_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_11[10] = dl_detect_out ? proc_dep_vld_vec_11_reg[10] : (proc_11_data_FIFO_blk[10] | proc_11_data_PIPO_blk[10] | proc_11_start_FIFO_blk[10] | proc_11_TLF_FIFO_blk[10] | proc_11_input_sync_blk[10] | proc_11_output_sync_blk[10]);
    assign proc_11_data_FIFO_blk[11] = 1'b0;
    assign proc_11_data_PIPO_blk[11] = 1'b0;
    assign proc_11_start_FIFO_blk[11] = 1'b0;
    assign proc_11_TLF_FIFO_blk[11] = 1'b0;
    assign proc_11_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_11_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_11[11] = dl_detect_out ? proc_dep_vld_vec_11_reg[11] : (proc_11_data_FIFO_blk[11] | proc_11_data_PIPO_blk[11] | proc_11_start_FIFO_blk[11] | proc_11_TLF_FIFO_blk[11] | proc_11_input_sync_blk[11] | proc_11_output_sync_blk[11]);
    assign proc_11_data_FIFO_blk[12] = 1'b0;
    assign proc_11_data_PIPO_blk[12] = 1'b0;
    assign proc_11_start_FIFO_blk[12] = 1'b0;
    assign proc_11_TLF_FIFO_blk[12] = 1'b0;
    assign proc_11_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_11_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_11[12] = dl_detect_out ? proc_dep_vld_vec_11_reg[12] : (proc_11_data_FIFO_blk[12] | proc_11_data_PIPO_blk[12] | proc_11_start_FIFO_blk[12] | proc_11_TLF_FIFO_blk[12] | proc_11_input_sync_blk[12] | proc_11_output_sync_blk[12]);
    assign proc_11_data_FIFO_blk[13] = 1'b0;
    assign proc_11_data_PIPO_blk[13] = 1'b0;
    assign proc_11_start_FIFO_blk[13] = 1'b0;
    assign proc_11_TLF_FIFO_blk[13] = 1'b0;
    assign proc_11_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_11_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_11[13] = dl_detect_out ? proc_dep_vld_vec_11_reg[13] : (proc_11_data_FIFO_blk[13] | proc_11_data_PIPO_blk[13] | proc_11_start_FIFO_blk[13] | proc_11_TLF_FIFO_blk[13] | proc_11_input_sync_blk[13] | proc_11_output_sync_blk[13]);
    assign proc_11_data_FIFO_blk[14] = 1'b0;
    assign proc_11_data_PIPO_blk[14] = 1'b0;
    assign proc_11_start_FIFO_blk[14] = 1'b0;
    assign proc_11_TLF_FIFO_blk[14] = 1'b0;
    assign proc_11_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_11_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_11[14] = dl_detect_out ? proc_dep_vld_vec_11_reg[14] : (proc_11_data_FIFO_blk[14] | proc_11_data_PIPO_blk[14] | proc_11_start_FIFO_blk[14] | proc_11_TLF_FIFO_blk[14] | proc_11_input_sync_blk[14] | proc_11_output_sync_blk[14]);
    assign proc_11_data_FIFO_blk[15] = 1'b0;
    assign proc_11_data_PIPO_blk[15] = 1'b0;
    assign proc_11_start_FIFO_blk[15] = 1'b0;
    assign proc_11_TLF_FIFO_blk[15] = 1'b0;
    assign proc_11_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_11_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_11[15] = dl_detect_out ? proc_dep_vld_vec_11_reg[15] : (proc_11_data_FIFO_blk[15] | proc_11_data_PIPO_blk[15] | proc_11_start_FIFO_blk[15] | proc_11_TLF_FIFO_blk[15] | proc_11_input_sync_blk[15] | proc_11_output_sync_blk[15]);
    assign proc_11_data_FIFO_blk[16] = 1'b0;
    assign proc_11_data_PIPO_blk[16] = 1'b0;
    assign proc_11_start_FIFO_blk[16] = 1'b0;
    assign proc_11_TLF_FIFO_blk[16] = 1'b0;
    assign proc_11_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_11_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_11[16] = dl_detect_out ? proc_dep_vld_vec_11_reg[16] : (proc_11_data_FIFO_blk[16] | proc_11_data_PIPO_blk[16] | proc_11_start_FIFO_blk[16] | proc_11_TLF_FIFO_blk[16] | proc_11_input_sync_blk[16] | proc_11_output_sync_blk[16]);
    assign proc_11_data_FIFO_blk[17] = 1'b0;
    assign proc_11_data_PIPO_blk[17] = 1'b0;
    assign proc_11_start_FIFO_blk[17] = 1'b0;
    assign proc_11_TLF_FIFO_blk[17] = 1'b0;
    assign proc_11_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_11_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_11[17] = dl_detect_out ? proc_dep_vld_vec_11_reg[17] : (proc_11_data_FIFO_blk[17] | proc_11_data_PIPO_blk[17] | proc_11_start_FIFO_blk[17] | proc_11_TLF_FIFO_blk[17] | proc_11_input_sync_blk[17] | proc_11_output_sync_blk[17]);
    assign proc_11_data_FIFO_blk[18] = 1'b0;
    assign proc_11_data_PIPO_blk[18] = 1'b0;
    assign proc_11_start_FIFO_blk[18] = 1'b0;
    assign proc_11_TLF_FIFO_blk[18] = 1'b0;
    assign proc_11_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_11_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_11[18] = dl_detect_out ? proc_dep_vld_vec_11_reg[18] : (proc_11_data_FIFO_blk[18] | proc_11_data_PIPO_blk[18] | proc_11_start_FIFO_blk[18] | proc_11_TLF_FIFO_blk[18] | proc_11_input_sync_blk[18] | proc_11_output_sync_blk[18]);
    assign proc_11_data_FIFO_blk[19] = 1'b0;
    assign proc_11_data_PIPO_blk[19] = 1'b0;
    assign proc_11_start_FIFO_blk[19] = 1'b0;
    assign proc_11_TLF_FIFO_blk[19] = 1'b0;
    assign proc_11_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_11_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_11[19] = dl_detect_out ? proc_dep_vld_vec_11_reg[19] : (proc_11_data_FIFO_blk[19] | proc_11_data_PIPO_blk[19] | proc_11_start_FIFO_blk[19] | proc_11_TLF_FIFO_blk[19] | proc_11_input_sync_blk[19] | proc_11_output_sync_blk[19]);
    assign proc_11_data_FIFO_blk[20] = 1'b0;
    assign proc_11_data_PIPO_blk[20] = 1'b0;
    assign proc_11_start_FIFO_blk[20] = 1'b0;
    assign proc_11_TLF_FIFO_blk[20] = 1'b0;
    assign proc_11_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_11_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_11[20] = dl_detect_out ? proc_dep_vld_vec_11_reg[20] : (proc_11_data_FIFO_blk[20] | proc_11_data_PIPO_blk[20] | proc_11_start_FIFO_blk[20] | proc_11_TLF_FIFO_blk[20] | proc_11_input_sync_blk[20] | proc_11_output_sync_blk[20]);
    assign proc_11_data_FIFO_blk[21] = 1'b0;
    assign proc_11_data_PIPO_blk[21] = 1'b0;
    assign proc_11_start_FIFO_blk[21] = 1'b0;
    assign proc_11_TLF_FIFO_blk[21] = 1'b0;
    assign proc_11_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_11_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_11[21] = dl_detect_out ? proc_dep_vld_vec_11_reg[21] : (proc_11_data_FIFO_blk[21] | proc_11_data_PIPO_blk[21] | proc_11_start_FIFO_blk[21] | proc_11_TLF_FIFO_blk[21] | proc_11_input_sync_blk[21] | proc_11_output_sync_blk[21]);
    assign proc_11_data_FIFO_blk[22] = 1'b0;
    assign proc_11_data_PIPO_blk[22] = 1'b0;
    assign proc_11_start_FIFO_blk[22] = 1'b0;
    assign proc_11_TLF_FIFO_blk[22] = 1'b0;
    assign proc_11_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_11_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_11[22] = dl_detect_out ? proc_dep_vld_vec_11_reg[22] : (proc_11_data_FIFO_blk[22] | proc_11_data_PIPO_blk[22] | proc_11_start_FIFO_blk[22] | proc_11_TLF_FIFO_blk[22] | proc_11_input_sync_blk[22] | proc_11_output_sync_blk[22]);
    assign proc_11_data_FIFO_blk[23] = 1'b0;
    assign proc_11_data_PIPO_blk[23] = 1'b0;
    assign proc_11_start_FIFO_blk[23] = 1'b0;
    assign proc_11_TLF_FIFO_blk[23] = 1'b0;
    assign proc_11_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_11_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_11[23] = dl_detect_out ? proc_dep_vld_vec_11_reg[23] : (proc_11_data_FIFO_blk[23] | proc_11_data_PIPO_blk[23] | proc_11_start_FIFO_blk[23] | proc_11_TLF_FIFO_blk[23] | proc_11_input_sync_blk[23] | proc_11_output_sync_blk[23]);
    assign proc_11_data_FIFO_blk[24] = 1'b0;
    assign proc_11_data_PIPO_blk[24] = 1'b0;
    assign proc_11_start_FIFO_blk[24] = 1'b0;
    assign proc_11_TLF_FIFO_blk[24] = 1'b0;
    assign proc_11_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_11_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_11[24] = dl_detect_out ? proc_dep_vld_vec_11_reg[24] : (proc_11_data_FIFO_blk[24] | proc_11_data_PIPO_blk[24] | proc_11_start_FIFO_blk[24] | proc_11_TLF_FIFO_blk[24] | proc_11_input_sync_blk[24] | proc_11_output_sync_blk[24]);
    assign proc_11_data_FIFO_blk[25] = 1'b0;
    assign proc_11_data_PIPO_blk[25] = 1'b0;
    assign proc_11_start_FIFO_blk[25] = 1'b0;
    assign proc_11_TLF_FIFO_blk[25] = 1'b0;
    assign proc_11_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_11_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_11[25] = dl_detect_out ? proc_dep_vld_vec_11_reg[25] : (proc_11_data_FIFO_blk[25] | proc_11_data_PIPO_blk[25] | proc_11_start_FIFO_blk[25] | proc_11_TLF_FIFO_blk[25] | proc_11_input_sync_blk[25] | proc_11_output_sync_blk[25]);
    assign proc_11_data_FIFO_blk[26] = 1'b0;
    assign proc_11_data_PIPO_blk[26] = 1'b0;
    assign proc_11_start_FIFO_blk[26] = 1'b0;
    assign proc_11_TLF_FIFO_blk[26] = 1'b0;
    assign proc_11_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_11_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_11[26] = dl_detect_out ? proc_dep_vld_vec_11_reg[26] : (proc_11_data_FIFO_blk[26] | proc_11_data_PIPO_blk[26] | proc_11_start_FIFO_blk[26] | proc_11_TLF_FIFO_blk[26] | proc_11_input_sync_blk[26] | proc_11_output_sync_blk[26]);
    assign proc_11_data_FIFO_blk[27] = 1'b0;
    assign proc_11_data_PIPO_blk[27] = 1'b0;
    assign proc_11_start_FIFO_blk[27] = 1'b0;
    assign proc_11_TLF_FIFO_blk[27] = 1'b0;
    assign proc_11_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_11_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_11[27] = dl_detect_out ? proc_dep_vld_vec_11_reg[27] : (proc_11_data_FIFO_blk[27] | proc_11_data_PIPO_blk[27] | proc_11_start_FIFO_blk[27] | proc_11_TLF_FIFO_blk[27] | proc_11_input_sync_blk[27] | proc_11_output_sync_blk[27]);
    assign proc_11_data_FIFO_blk[28] = 1'b0;
    assign proc_11_data_PIPO_blk[28] = 1'b0;
    assign proc_11_start_FIFO_blk[28] = 1'b0;
    assign proc_11_TLF_FIFO_blk[28] = 1'b0;
    assign proc_11_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_11_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_11[28] = dl_detect_out ? proc_dep_vld_vec_11_reg[28] : (proc_11_data_FIFO_blk[28] | proc_11_data_PIPO_blk[28] | proc_11_start_FIFO_blk[28] | proc_11_TLF_FIFO_blk[28] | proc_11_input_sync_blk[28] | proc_11_output_sync_blk[28]);
    assign proc_11_data_FIFO_blk[29] = 1'b0;
    assign proc_11_data_PIPO_blk[29] = 1'b0;
    assign proc_11_start_FIFO_blk[29] = 1'b0;
    assign proc_11_TLF_FIFO_blk[29] = 1'b0;
    assign proc_11_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_11_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_11[29] = dl_detect_out ? proc_dep_vld_vec_11_reg[29] : (proc_11_data_FIFO_blk[29] | proc_11_data_PIPO_blk[29] | proc_11_start_FIFO_blk[29] | proc_11_TLF_FIFO_blk[29] | proc_11_input_sync_blk[29] | proc_11_output_sync_blk[29]);
    assign proc_11_data_FIFO_blk[30] = 1'b0;
    assign proc_11_data_PIPO_blk[30] = 1'b0;
    assign proc_11_start_FIFO_blk[30] = 1'b0;
    assign proc_11_TLF_FIFO_blk[30] = 1'b0;
    assign proc_11_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_11_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_11[30] = dl_detect_out ? proc_dep_vld_vec_11_reg[30] : (proc_11_data_FIFO_blk[30] | proc_11_data_PIPO_blk[30] | proc_11_start_FIFO_blk[30] | proc_11_TLF_FIFO_blk[30] | proc_11_input_sync_blk[30] | proc_11_output_sync_blk[30]);
    assign proc_11_data_FIFO_blk[31] = 1'b0;
    assign proc_11_data_PIPO_blk[31] = 1'b0;
    assign proc_11_start_FIFO_blk[31] = 1'b0;
    assign proc_11_TLF_FIFO_blk[31] = 1'b0;
    assign proc_11_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_11_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_11[31] = dl_detect_out ? proc_dep_vld_vec_11_reg[31] : (proc_11_data_FIFO_blk[31] | proc_11_data_PIPO_blk[31] | proc_11_start_FIFO_blk[31] | proc_11_TLF_FIFO_blk[31] | proc_11_input_sync_blk[31] | proc_11_output_sync_blk[31]);
    assign proc_11_data_FIFO_blk[32] = 1'b0;
    assign proc_11_data_PIPO_blk[32] = 1'b0;
    assign proc_11_start_FIFO_blk[32] = 1'b0;
    assign proc_11_TLF_FIFO_blk[32] = 1'b0;
    assign proc_11_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_6_U0_ap_ready & ProcessingElement_6_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_11_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_11[32] = dl_detect_out ? proc_dep_vld_vec_11_reg[32] : (proc_11_data_FIFO_blk[32] | proc_11_data_PIPO_blk[32] | proc_11_start_FIFO_blk[32] | proc_11_TLF_FIFO_blk[32] | proc_11_input_sync_blk[32] | proc_11_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_11_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_11_reg <= proc_dep_vld_vec_11;
        end
    end
    assign in_chan_dep_vld_vec_11[0] = dep_chan_vld_0_11;
    assign in_chan_dep_data_vec_11[39 : 0] = dep_chan_data_0_11;
    assign token_in_vec_11[0] = token_0_11;
    assign in_chan_dep_vld_vec_11[1] = dep_chan_vld_1_11;
    assign in_chan_dep_data_vec_11[79 : 40] = dep_chan_data_1_11;
    assign token_in_vec_11[1] = token_1_11;
    assign in_chan_dep_vld_vec_11[2] = dep_chan_vld_3_11;
    assign in_chan_dep_data_vec_11[119 : 80] = dep_chan_data_3_11;
    assign token_in_vec_11[2] = token_3_11;
    assign in_chan_dep_vld_vec_11[3] = dep_chan_vld_6_11;
    assign in_chan_dep_data_vec_11[159 : 120] = dep_chan_data_6_11;
    assign token_in_vec_11[3] = token_6_11;
    assign in_chan_dep_vld_vec_11[4] = dep_chan_vld_7_11;
    assign in_chan_dep_data_vec_11[199 : 160] = dep_chan_data_7_11;
    assign token_in_vec_11[4] = token_7_11;
    assign in_chan_dep_vld_vec_11[5] = dep_chan_vld_8_11;
    assign in_chan_dep_data_vec_11[239 : 200] = dep_chan_data_8_11;
    assign token_in_vec_11[5] = token_8_11;
    assign in_chan_dep_vld_vec_11[6] = dep_chan_vld_9_11;
    assign in_chan_dep_data_vec_11[279 : 240] = dep_chan_data_9_11;
    assign token_in_vec_11[6] = token_9_11;
    assign in_chan_dep_vld_vec_11[7] = dep_chan_vld_10_11;
    assign in_chan_dep_data_vec_11[319 : 280] = dep_chan_data_10_11;
    assign token_in_vec_11[7] = token_10_11;
    assign in_chan_dep_vld_vec_11[8] = dep_chan_vld_12_11;
    assign in_chan_dep_data_vec_11[359 : 320] = dep_chan_data_12_11;
    assign token_in_vec_11[8] = token_12_11;
    assign in_chan_dep_vld_vec_11[9] = dep_chan_vld_13_11;
    assign in_chan_dep_data_vec_11[399 : 360] = dep_chan_data_13_11;
    assign token_in_vec_11[9] = token_13_11;
    assign in_chan_dep_vld_vec_11[10] = dep_chan_vld_14_11;
    assign in_chan_dep_data_vec_11[439 : 400] = dep_chan_data_14_11;
    assign token_in_vec_11[10] = token_14_11;
    assign in_chan_dep_vld_vec_11[11] = dep_chan_vld_15_11;
    assign in_chan_dep_data_vec_11[479 : 440] = dep_chan_data_15_11;
    assign token_in_vec_11[11] = token_15_11;
    assign in_chan_dep_vld_vec_11[12] = dep_chan_vld_16_11;
    assign in_chan_dep_data_vec_11[519 : 480] = dep_chan_data_16_11;
    assign token_in_vec_11[12] = token_16_11;
    assign in_chan_dep_vld_vec_11[13] = dep_chan_vld_17_11;
    assign in_chan_dep_data_vec_11[559 : 520] = dep_chan_data_17_11;
    assign token_in_vec_11[13] = token_17_11;
    assign in_chan_dep_vld_vec_11[14] = dep_chan_vld_18_11;
    assign in_chan_dep_data_vec_11[599 : 560] = dep_chan_data_18_11;
    assign token_in_vec_11[14] = token_18_11;
    assign in_chan_dep_vld_vec_11[15] = dep_chan_vld_19_11;
    assign in_chan_dep_data_vec_11[639 : 600] = dep_chan_data_19_11;
    assign token_in_vec_11[15] = token_19_11;
    assign in_chan_dep_vld_vec_11[16] = dep_chan_vld_20_11;
    assign in_chan_dep_data_vec_11[679 : 640] = dep_chan_data_20_11;
    assign token_in_vec_11[16] = token_20_11;
    assign in_chan_dep_vld_vec_11[17] = dep_chan_vld_21_11;
    assign in_chan_dep_data_vec_11[719 : 680] = dep_chan_data_21_11;
    assign token_in_vec_11[17] = token_21_11;
    assign in_chan_dep_vld_vec_11[18] = dep_chan_vld_22_11;
    assign in_chan_dep_data_vec_11[759 : 720] = dep_chan_data_22_11;
    assign token_in_vec_11[18] = token_22_11;
    assign in_chan_dep_vld_vec_11[19] = dep_chan_vld_23_11;
    assign in_chan_dep_data_vec_11[799 : 760] = dep_chan_data_23_11;
    assign token_in_vec_11[19] = token_23_11;
    assign in_chan_dep_vld_vec_11[20] = dep_chan_vld_24_11;
    assign in_chan_dep_data_vec_11[839 : 800] = dep_chan_data_24_11;
    assign token_in_vec_11[20] = token_24_11;
    assign in_chan_dep_vld_vec_11[21] = dep_chan_vld_25_11;
    assign in_chan_dep_data_vec_11[879 : 840] = dep_chan_data_25_11;
    assign token_in_vec_11[21] = token_25_11;
    assign in_chan_dep_vld_vec_11[22] = dep_chan_vld_26_11;
    assign in_chan_dep_data_vec_11[919 : 880] = dep_chan_data_26_11;
    assign token_in_vec_11[22] = token_26_11;
    assign in_chan_dep_vld_vec_11[23] = dep_chan_vld_27_11;
    assign in_chan_dep_data_vec_11[959 : 920] = dep_chan_data_27_11;
    assign token_in_vec_11[23] = token_27_11;
    assign in_chan_dep_vld_vec_11[24] = dep_chan_vld_28_11;
    assign in_chan_dep_data_vec_11[999 : 960] = dep_chan_data_28_11;
    assign token_in_vec_11[24] = token_28_11;
    assign in_chan_dep_vld_vec_11[25] = dep_chan_vld_29_11;
    assign in_chan_dep_data_vec_11[1039 : 1000] = dep_chan_data_29_11;
    assign token_in_vec_11[25] = token_29_11;
    assign in_chan_dep_vld_vec_11[26] = dep_chan_vld_30_11;
    assign in_chan_dep_data_vec_11[1079 : 1040] = dep_chan_data_30_11;
    assign token_in_vec_11[26] = token_30_11;
    assign in_chan_dep_vld_vec_11[27] = dep_chan_vld_31_11;
    assign in_chan_dep_data_vec_11[1119 : 1080] = dep_chan_data_31_11;
    assign token_in_vec_11[27] = token_31_11;
    assign in_chan_dep_vld_vec_11[28] = dep_chan_vld_32_11;
    assign in_chan_dep_data_vec_11[1159 : 1120] = dep_chan_data_32_11;
    assign token_in_vec_11[28] = token_32_11;
    assign in_chan_dep_vld_vec_11[29] = dep_chan_vld_33_11;
    assign in_chan_dep_data_vec_11[1199 : 1160] = dep_chan_data_33_11;
    assign token_in_vec_11[29] = token_33_11;
    assign in_chan_dep_vld_vec_11[30] = dep_chan_vld_34_11;
    assign in_chan_dep_data_vec_11[1239 : 1200] = dep_chan_data_34_11;
    assign token_in_vec_11[30] = token_34_11;
    assign in_chan_dep_vld_vec_11[31] = dep_chan_vld_35_11;
    assign in_chan_dep_data_vec_11[1279 : 1240] = dep_chan_data_35_11;
    assign token_in_vec_11[31] = token_35_11;
    assign in_chan_dep_vld_vec_11[32] = dep_chan_vld_36_11;
    assign in_chan_dep_data_vec_11[1319 : 1280] = dep_chan_data_36_11;
    assign token_in_vec_11[32] = token_36_11;
    assign dep_chan_vld_11_10 = out_chan_dep_vld_vec_11[0];
    assign dep_chan_data_11_10 = out_chan_dep_data_11;
    assign token_11_10 = token_out_vec_11[0];
    assign dep_chan_vld_11_12 = out_chan_dep_vld_vec_11[1];
    assign dep_chan_data_11_12 = out_chan_dep_data_11;
    assign token_11_12 = token_out_vec_11[1];
    assign dep_chan_vld_11_0 = out_chan_dep_vld_vec_11[2];
    assign dep_chan_data_11_0 = out_chan_dep_data_11;
    assign token_11_0 = token_out_vec_11[2];
    assign dep_chan_vld_11_1 = out_chan_dep_vld_vec_11[3];
    assign dep_chan_data_11_1 = out_chan_dep_data_11;
    assign token_11_1 = token_out_vec_11[3];
    assign dep_chan_vld_11_3 = out_chan_dep_vld_vec_11[4];
    assign dep_chan_data_11_3 = out_chan_dep_data_11;
    assign token_11_3 = token_out_vec_11[4];
    assign dep_chan_vld_11_6 = out_chan_dep_vld_vec_11[5];
    assign dep_chan_data_11_6 = out_chan_dep_data_11;
    assign token_11_6 = token_out_vec_11[5];
    assign dep_chan_vld_11_7 = out_chan_dep_vld_vec_11[6];
    assign dep_chan_data_11_7 = out_chan_dep_data_11;
    assign token_11_7 = token_out_vec_11[6];
    assign dep_chan_vld_11_8 = out_chan_dep_vld_vec_11[7];
    assign dep_chan_data_11_8 = out_chan_dep_data_11;
    assign token_11_8 = token_out_vec_11[7];
    assign dep_chan_vld_11_9 = out_chan_dep_vld_vec_11[8];
    assign dep_chan_data_11_9 = out_chan_dep_data_11;
    assign token_11_9 = token_out_vec_11[8];
    assign dep_chan_vld_11_13 = out_chan_dep_vld_vec_11[9];
    assign dep_chan_data_11_13 = out_chan_dep_data_11;
    assign token_11_13 = token_out_vec_11[9];
    assign dep_chan_vld_11_14 = out_chan_dep_vld_vec_11[10];
    assign dep_chan_data_11_14 = out_chan_dep_data_11;
    assign token_11_14 = token_out_vec_11[10];
    assign dep_chan_vld_11_15 = out_chan_dep_vld_vec_11[11];
    assign dep_chan_data_11_15 = out_chan_dep_data_11;
    assign token_11_15 = token_out_vec_11[11];
    assign dep_chan_vld_11_16 = out_chan_dep_vld_vec_11[12];
    assign dep_chan_data_11_16 = out_chan_dep_data_11;
    assign token_11_16 = token_out_vec_11[12];
    assign dep_chan_vld_11_17 = out_chan_dep_vld_vec_11[13];
    assign dep_chan_data_11_17 = out_chan_dep_data_11;
    assign token_11_17 = token_out_vec_11[13];
    assign dep_chan_vld_11_18 = out_chan_dep_vld_vec_11[14];
    assign dep_chan_data_11_18 = out_chan_dep_data_11;
    assign token_11_18 = token_out_vec_11[14];
    assign dep_chan_vld_11_19 = out_chan_dep_vld_vec_11[15];
    assign dep_chan_data_11_19 = out_chan_dep_data_11;
    assign token_11_19 = token_out_vec_11[15];
    assign dep_chan_vld_11_20 = out_chan_dep_vld_vec_11[16];
    assign dep_chan_data_11_20 = out_chan_dep_data_11;
    assign token_11_20 = token_out_vec_11[16];
    assign dep_chan_vld_11_21 = out_chan_dep_vld_vec_11[17];
    assign dep_chan_data_11_21 = out_chan_dep_data_11;
    assign token_11_21 = token_out_vec_11[17];
    assign dep_chan_vld_11_22 = out_chan_dep_vld_vec_11[18];
    assign dep_chan_data_11_22 = out_chan_dep_data_11;
    assign token_11_22 = token_out_vec_11[18];
    assign dep_chan_vld_11_23 = out_chan_dep_vld_vec_11[19];
    assign dep_chan_data_11_23 = out_chan_dep_data_11;
    assign token_11_23 = token_out_vec_11[19];
    assign dep_chan_vld_11_24 = out_chan_dep_vld_vec_11[20];
    assign dep_chan_data_11_24 = out_chan_dep_data_11;
    assign token_11_24 = token_out_vec_11[20];
    assign dep_chan_vld_11_25 = out_chan_dep_vld_vec_11[21];
    assign dep_chan_data_11_25 = out_chan_dep_data_11;
    assign token_11_25 = token_out_vec_11[21];
    assign dep_chan_vld_11_26 = out_chan_dep_vld_vec_11[22];
    assign dep_chan_data_11_26 = out_chan_dep_data_11;
    assign token_11_26 = token_out_vec_11[22];
    assign dep_chan_vld_11_27 = out_chan_dep_vld_vec_11[23];
    assign dep_chan_data_11_27 = out_chan_dep_data_11;
    assign token_11_27 = token_out_vec_11[23];
    assign dep_chan_vld_11_28 = out_chan_dep_vld_vec_11[24];
    assign dep_chan_data_11_28 = out_chan_dep_data_11;
    assign token_11_28 = token_out_vec_11[24];
    assign dep_chan_vld_11_29 = out_chan_dep_vld_vec_11[25];
    assign dep_chan_data_11_29 = out_chan_dep_data_11;
    assign token_11_29 = token_out_vec_11[25];
    assign dep_chan_vld_11_30 = out_chan_dep_vld_vec_11[26];
    assign dep_chan_data_11_30 = out_chan_dep_data_11;
    assign token_11_30 = token_out_vec_11[26];
    assign dep_chan_vld_11_31 = out_chan_dep_vld_vec_11[27];
    assign dep_chan_data_11_31 = out_chan_dep_data_11;
    assign token_11_31 = token_out_vec_11[27];
    assign dep_chan_vld_11_32 = out_chan_dep_vld_vec_11[28];
    assign dep_chan_data_11_32 = out_chan_dep_data_11;
    assign token_11_32 = token_out_vec_11[28];
    assign dep_chan_vld_11_33 = out_chan_dep_vld_vec_11[29];
    assign dep_chan_data_11_33 = out_chan_dep_data_11;
    assign token_11_33 = token_out_vec_11[29];
    assign dep_chan_vld_11_34 = out_chan_dep_vld_vec_11[30];
    assign dep_chan_data_11_34 = out_chan_dep_data_11;
    assign token_11_34 = token_out_vec_11[30];
    assign dep_chan_vld_11_35 = out_chan_dep_vld_vec_11[31];
    assign dep_chan_data_11_35 = out_chan_dep_data_11;
    assign token_11_35 = token_out_vec_11[31];
    assign dep_chan_vld_11_36 = out_chan_dep_vld_vec_11[32];
    assign dep_chan_data_11_36 = out_chan_dep_data_11;
    assign token_11_36 = token_out_vec_11[32];

    // Process: ProcessingElement_7_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 12, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_12 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_12),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_12),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_12),
        .token_in_vec(token_in_vec_12),
        .dl_detect_in(dl_detect_out),
        .origin(origin[12]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_12),
        .out_chan_dep_data(out_chan_dep_data_12),
        .token_out_vec(token_out_vec_12),
        .dl_detect_out(dl_in_vec[12]));

    assign proc_12_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_6_blk_n) | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_6_blk_n) | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_WriteC_Flattened_fu_179.cPipes_6_blk_n);
    assign proc_12_data_PIPO_blk[0] = 1'b0;
    assign proc_12_start_FIFO_blk[0] = 1'b0;
    assign proc_12_TLF_FIFO_blk[0] = 1'b0;
    assign proc_12_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_12_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_12[0] = dl_detect_out ? proc_dep_vld_vec_12_reg[0] : (proc_12_data_FIFO_blk[0] | proc_12_data_PIPO_blk[0] | proc_12_start_FIFO_blk[0] | proc_12_TLF_FIFO_blk[0] | proc_12_input_sync_blk[0] | proc_12_output_sync_blk[0]);
    assign proc_12_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_7_blk_n) | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_7_blk_n) | (~ProcessingElement_7_U0.grp_ProcessingElement_7_Pipeline_WriteC_Flattened_fu_179.cPipes_7_blk_n);
    assign proc_12_data_PIPO_blk[1] = 1'b0;
    assign proc_12_start_FIFO_blk[1] = 1'b0;
    assign proc_12_TLF_FIFO_blk[1] = 1'b0;
    assign proc_12_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_12_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_12[1] = dl_detect_out ? proc_dep_vld_vec_12_reg[1] : (proc_12_data_FIFO_blk[1] | proc_12_data_PIPO_blk[1] | proc_12_start_FIFO_blk[1] | proc_12_TLF_FIFO_blk[1] | proc_12_input_sync_blk[1] | proc_12_output_sync_blk[1]);
    assign proc_12_data_FIFO_blk[2] = 1'b0;
    assign proc_12_data_PIPO_blk[2] = 1'b0;
    assign proc_12_start_FIFO_blk[2] = 1'b0;
    assign proc_12_TLF_FIFO_blk[2] = 1'b0;
    assign proc_12_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_12_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_12[2] = dl_detect_out ? proc_dep_vld_vec_12_reg[2] : (proc_12_data_FIFO_blk[2] | proc_12_data_PIPO_blk[2] | proc_12_start_FIFO_blk[2] | proc_12_TLF_FIFO_blk[2] | proc_12_input_sync_blk[2] | proc_12_output_sync_blk[2]);
    assign proc_12_data_FIFO_blk[3] = 1'b0;
    assign proc_12_data_PIPO_blk[3] = 1'b0;
    assign proc_12_start_FIFO_blk[3] = 1'b0;
    assign proc_12_TLF_FIFO_blk[3] = 1'b0;
    assign proc_12_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_12_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_12[3] = dl_detect_out ? proc_dep_vld_vec_12_reg[3] : (proc_12_data_FIFO_blk[3] | proc_12_data_PIPO_blk[3] | proc_12_start_FIFO_blk[3] | proc_12_TLF_FIFO_blk[3] | proc_12_input_sync_blk[3] | proc_12_output_sync_blk[3]);
    assign proc_12_data_FIFO_blk[4] = 1'b0;
    assign proc_12_data_PIPO_blk[4] = 1'b0;
    assign proc_12_start_FIFO_blk[4] = 1'b0;
    assign proc_12_TLF_FIFO_blk[4] = 1'b0;
    assign proc_12_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_12_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_12[4] = dl_detect_out ? proc_dep_vld_vec_12_reg[4] : (proc_12_data_FIFO_blk[4] | proc_12_data_PIPO_blk[4] | proc_12_start_FIFO_blk[4] | proc_12_TLF_FIFO_blk[4] | proc_12_input_sync_blk[4] | proc_12_output_sync_blk[4]);
    assign proc_12_data_FIFO_blk[5] = 1'b0;
    assign proc_12_data_PIPO_blk[5] = 1'b0;
    assign proc_12_start_FIFO_blk[5] = 1'b0;
    assign proc_12_TLF_FIFO_blk[5] = 1'b0;
    assign proc_12_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_12_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_12[5] = dl_detect_out ? proc_dep_vld_vec_12_reg[5] : (proc_12_data_FIFO_blk[5] | proc_12_data_PIPO_blk[5] | proc_12_start_FIFO_blk[5] | proc_12_TLF_FIFO_blk[5] | proc_12_input_sync_blk[5] | proc_12_output_sync_blk[5]);
    assign proc_12_data_FIFO_blk[6] = 1'b0;
    assign proc_12_data_PIPO_blk[6] = 1'b0;
    assign proc_12_start_FIFO_blk[6] = 1'b0;
    assign proc_12_TLF_FIFO_blk[6] = 1'b0;
    assign proc_12_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_12_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_12[6] = dl_detect_out ? proc_dep_vld_vec_12_reg[6] : (proc_12_data_FIFO_blk[6] | proc_12_data_PIPO_blk[6] | proc_12_start_FIFO_blk[6] | proc_12_TLF_FIFO_blk[6] | proc_12_input_sync_blk[6] | proc_12_output_sync_blk[6]);
    assign proc_12_data_FIFO_blk[7] = 1'b0;
    assign proc_12_data_PIPO_blk[7] = 1'b0;
    assign proc_12_start_FIFO_blk[7] = 1'b0;
    assign proc_12_TLF_FIFO_blk[7] = 1'b0;
    assign proc_12_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_12_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_12[7] = dl_detect_out ? proc_dep_vld_vec_12_reg[7] : (proc_12_data_FIFO_blk[7] | proc_12_data_PIPO_blk[7] | proc_12_start_FIFO_blk[7] | proc_12_TLF_FIFO_blk[7] | proc_12_input_sync_blk[7] | proc_12_output_sync_blk[7]);
    assign proc_12_data_FIFO_blk[8] = 1'b0;
    assign proc_12_data_PIPO_blk[8] = 1'b0;
    assign proc_12_start_FIFO_blk[8] = 1'b0;
    assign proc_12_TLF_FIFO_blk[8] = 1'b0;
    assign proc_12_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_12_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_12[8] = dl_detect_out ? proc_dep_vld_vec_12_reg[8] : (proc_12_data_FIFO_blk[8] | proc_12_data_PIPO_blk[8] | proc_12_start_FIFO_blk[8] | proc_12_TLF_FIFO_blk[8] | proc_12_input_sync_blk[8] | proc_12_output_sync_blk[8]);
    assign proc_12_data_FIFO_blk[9] = 1'b0;
    assign proc_12_data_PIPO_blk[9] = 1'b0;
    assign proc_12_start_FIFO_blk[9] = 1'b0;
    assign proc_12_TLF_FIFO_blk[9] = 1'b0;
    assign proc_12_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_12_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_12[9] = dl_detect_out ? proc_dep_vld_vec_12_reg[9] : (proc_12_data_FIFO_blk[9] | proc_12_data_PIPO_blk[9] | proc_12_start_FIFO_blk[9] | proc_12_TLF_FIFO_blk[9] | proc_12_input_sync_blk[9] | proc_12_output_sync_blk[9]);
    assign proc_12_data_FIFO_blk[10] = 1'b0;
    assign proc_12_data_PIPO_blk[10] = 1'b0;
    assign proc_12_start_FIFO_blk[10] = 1'b0;
    assign proc_12_TLF_FIFO_blk[10] = 1'b0;
    assign proc_12_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_12_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_12[10] = dl_detect_out ? proc_dep_vld_vec_12_reg[10] : (proc_12_data_FIFO_blk[10] | proc_12_data_PIPO_blk[10] | proc_12_start_FIFO_blk[10] | proc_12_TLF_FIFO_blk[10] | proc_12_input_sync_blk[10] | proc_12_output_sync_blk[10]);
    assign proc_12_data_FIFO_blk[11] = 1'b0;
    assign proc_12_data_PIPO_blk[11] = 1'b0;
    assign proc_12_start_FIFO_blk[11] = 1'b0;
    assign proc_12_TLF_FIFO_blk[11] = 1'b0;
    assign proc_12_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_12_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_12[11] = dl_detect_out ? proc_dep_vld_vec_12_reg[11] : (proc_12_data_FIFO_blk[11] | proc_12_data_PIPO_blk[11] | proc_12_start_FIFO_blk[11] | proc_12_TLF_FIFO_blk[11] | proc_12_input_sync_blk[11] | proc_12_output_sync_blk[11]);
    assign proc_12_data_FIFO_blk[12] = 1'b0;
    assign proc_12_data_PIPO_blk[12] = 1'b0;
    assign proc_12_start_FIFO_blk[12] = 1'b0;
    assign proc_12_TLF_FIFO_blk[12] = 1'b0;
    assign proc_12_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_12_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_12[12] = dl_detect_out ? proc_dep_vld_vec_12_reg[12] : (proc_12_data_FIFO_blk[12] | proc_12_data_PIPO_blk[12] | proc_12_start_FIFO_blk[12] | proc_12_TLF_FIFO_blk[12] | proc_12_input_sync_blk[12] | proc_12_output_sync_blk[12]);
    assign proc_12_data_FIFO_blk[13] = 1'b0;
    assign proc_12_data_PIPO_blk[13] = 1'b0;
    assign proc_12_start_FIFO_blk[13] = 1'b0;
    assign proc_12_TLF_FIFO_blk[13] = 1'b0;
    assign proc_12_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_12_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_12[13] = dl_detect_out ? proc_dep_vld_vec_12_reg[13] : (proc_12_data_FIFO_blk[13] | proc_12_data_PIPO_blk[13] | proc_12_start_FIFO_blk[13] | proc_12_TLF_FIFO_blk[13] | proc_12_input_sync_blk[13] | proc_12_output_sync_blk[13]);
    assign proc_12_data_FIFO_blk[14] = 1'b0;
    assign proc_12_data_PIPO_blk[14] = 1'b0;
    assign proc_12_start_FIFO_blk[14] = 1'b0;
    assign proc_12_TLF_FIFO_blk[14] = 1'b0;
    assign proc_12_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_12_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_12[14] = dl_detect_out ? proc_dep_vld_vec_12_reg[14] : (proc_12_data_FIFO_blk[14] | proc_12_data_PIPO_blk[14] | proc_12_start_FIFO_blk[14] | proc_12_TLF_FIFO_blk[14] | proc_12_input_sync_blk[14] | proc_12_output_sync_blk[14]);
    assign proc_12_data_FIFO_blk[15] = 1'b0;
    assign proc_12_data_PIPO_blk[15] = 1'b0;
    assign proc_12_start_FIFO_blk[15] = 1'b0;
    assign proc_12_TLF_FIFO_blk[15] = 1'b0;
    assign proc_12_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_12_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_12[15] = dl_detect_out ? proc_dep_vld_vec_12_reg[15] : (proc_12_data_FIFO_blk[15] | proc_12_data_PIPO_blk[15] | proc_12_start_FIFO_blk[15] | proc_12_TLF_FIFO_blk[15] | proc_12_input_sync_blk[15] | proc_12_output_sync_blk[15]);
    assign proc_12_data_FIFO_blk[16] = 1'b0;
    assign proc_12_data_PIPO_blk[16] = 1'b0;
    assign proc_12_start_FIFO_blk[16] = 1'b0;
    assign proc_12_TLF_FIFO_blk[16] = 1'b0;
    assign proc_12_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_12_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_12[16] = dl_detect_out ? proc_dep_vld_vec_12_reg[16] : (proc_12_data_FIFO_blk[16] | proc_12_data_PIPO_blk[16] | proc_12_start_FIFO_blk[16] | proc_12_TLF_FIFO_blk[16] | proc_12_input_sync_blk[16] | proc_12_output_sync_blk[16]);
    assign proc_12_data_FIFO_blk[17] = 1'b0;
    assign proc_12_data_PIPO_blk[17] = 1'b0;
    assign proc_12_start_FIFO_blk[17] = 1'b0;
    assign proc_12_TLF_FIFO_blk[17] = 1'b0;
    assign proc_12_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_12_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_12[17] = dl_detect_out ? proc_dep_vld_vec_12_reg[17] : (proc_12_data_FIFO_blk[17] | proc_12_data_PIPO_blk[17] | proc_12_start_FIFO_blk[17] | proc_12_TLF_FIFO_blk[17] | proc_12_input_sync_blk[17] | proc_12_output_sync_blk[17]);
    assign proc_12_data_FIFO_blk[18] = 1'b0;
    assign proc_12_data_PIPO_blk[18] = 1'b0;
    assign proc_12_start_FIFO_blk[18] = 1'b0;
    assign proc_12_TLF_FIFO_blk[18] = 1'b0;
    assign proc_12_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_12_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_12[18] = dl_detect_out ? proc_dep_vld_vec_12_reg[18] : (proc_12_data_FIFO_blk[18] | proc_12_data_PIPO_blk[18] | proc_12_start_FIFO_blk[18] | proc_12_TLF_FIFO_blk[18] | proc_12_input_sync_blk[18] | proc_12_output_sync_blk[18]);
    assign proc_12_data_FIFO_blk[19] = 1'b0;
    assign proc_12_data_PIPO_blk[19] = 1'b0;
    assign proc_12_start_FIFO_blk[19] = 1'b0;
    assign proc_12_TLF_FIFO_blk[19] = 1'b0;
    assign proc_12_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_12_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_12[19] = dl_detect_out ? proc_dep_vld_vec_12_reg[19] : (proc_12_data_FIFO_blk[19] | proc_12_data_PIPO_blk[19] | proc_12_start_FIFO_blk[19] | proc_12_TLF_FIFO_blk[19] | proc_12_input_sync_blk[19] | proc_12_output_sync_blk[19]);
    assign proc_12_data_FIFO_blk[20] = 1'b0;
    assign proc_12_data_PIPO_blk[20] = 1'b0;
    assign proc_12_start_FIFO_blk[20] = 1'b0;
    assign proc_12_TLF_FIFO_blk[20] = 1'b0;
    assign proc_12_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_12_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_12[20] = dl_detect_out ? proc_dep_vld_vec_12_reg[20] : (proc_12_data_FIFO_blk[20] | proc_12_data_PIPO_blk[20] | proc_12_start_FIFO_blk[20] | proc_12_TLF_FIFO_blk[20] | proc_12_input_sync_blk[20] | proc_12_output_sync_blk[20]);
    assign proc_12_data_FIFO_blk[21] = 1'b0;
    assign proc_12_data_PIPO_blk[21] = 1'b0;
    assign proc_12_start_FIFO_blk[21] = 1'b0;
    assign proc_12_TLF_FIFO_blk[21] = 1'b0;
    assign proc_12_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_12_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_12[21] = dl_detect_out ? proc_dep_vld_vec_12_reg[21] : (proc_12_data_FIFO_blk[21] | proc_12_data_PIPO_blk[21] | proc_12_start_FIFO_blk[21] | proc_12_TLF_FIFO_blk[21] | proc_12_input_sync_blk[21] | proc_12_output_sync_blk[21]);
    assign proc_12_data_FIFO_blk[22] = 1'b0;
    assign proc_12_data_PIPO_blk[22] = 1'b0;
    assign proc_12_start_FIFO_blk[22] = 1'b0;
    assign proc_12_TLF_FIFO_blk[22] = 1'b0;
    assign proc_12_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_12_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_12[22] = dl_detect_out ? proc_dep_vld_vec_12_reg[22] : (proc_12_data_FIFO_blk[22] | proc_12_data_PIPO_blk[22] | proc_12_start_FIFO_blk[22] | proc_12_TLF_FIFO_blk[22] | proc_12_input_sync_blk[22] | proc_12_output_sync_blk[22]);
    assign proc_12_data_FIFO_blk[23] = 1'b0;
    assign proc_12_data_PIPO_blk[23] = 1'b0;
    assign proc_12_start_FIFO_blk[23] = 1'b0;
    assign proc_12_TLF_FIFO_blk[23] = 1'b0;
    assign proc_12_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_12_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_12[23] = dl_detect_out ? proc_dep_vld_vec_12_reg[23] : (proc_12_data_FIFO_blk[23] | proc_12_data_PIPO_blk[23] | proc_12_start_FIFO_blk[23] | proc_12_TLF_FIFO_blk[23] | proc_12_input_sync_blk[23] | proc_12_output_sync_blk[23]);
    assign proc_12_data_FIFO_blk[24] = 1'b0;
    assign proc_12_data_PIPO_blk[24] = 1'b0;
    assign proc_12_start_FIFO_blk[24] = 1'b0;
    assign proc_12_TLF_FIFO_blk[24] = 1'b0;
    assign proc_12_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_12_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_12[24] = dl_detect_out ? proc_dep_vld_vec_12_reg[24] : (proc_12_data_FIFO_blk[24] | proc_12_data_PIPO_blk[24] | proc_12_start_FIFO_blk[24] | proc_12_TLF_FIFO_blk[24] | proc_12_input_sync_blk[24] | proc_12_output_sync_blk[24]);
    assign proc_12_data_FIFO_blk[25] = 1'b0;
    assign proc_12_data_PIPO_blk[25] = 1'b0;
    assign proc_12_start_FIFO_blk[25] = 1'b0;
    assign proc_12_TLF_FIFO_blk[25] = 1'b0;
    assign proc_12_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_12_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_12[25] = dl_detect_out ? proc_dep_vld_vec_12_reg[25] : (proc_12_data_FIFO_blk[25] | proc_12_data_PIPO_blk[25] | proc_12_start_FIFO_blk[25] | proc_12_TLF_FIFO_blk[25] | proc_12_input_sync_blk[25] | proc_12_output_sync_blk[25]);
    assign proc_12_data_FIFO_blk[26] = 1'b0;
    assign proc_12_data_PIPO_blk[26] = 1'b0;
    assign proc_12_start_FIFO_blk[26] = 1'b0;
    assign proc_12_TLF_FIFO_blk[26] = 1'b0;
    assign proc_12_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_12_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_12[26] = dl_detect_out ? proc_dep_vld_vec_12_reg[26] : (proc_12_data_FIFO_blk[26] | proc_12_data_PIPO_blk[26] | proc_12_start_FIFO_blk[26] | proc_12_TLF_FIFO_blk[26] | proc_12_input_sync_blk[26] | proc_12_output_sync_blk[26]);
    assign proc_12_data_FIFO_blk[27] = 1'b0;
    assign proc_12_data_PIPO_blk[27] = 1'b0;
    assign proc_12_start_FIFO_blk[27] = 1'b0;
    assign proc_12_TLF_FIFO_blk[27] = 1'b0;
    assign proc_12_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_12_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_12[27] = dl_detect_out ? proc_dep_vld_vec_12_reg[27] : (proc_12_data_FIFO_blk[27] | proc_12_data_PIPO_blk[27] | proc_12_start_FIFO_blk[27] | proc_12_TLF_FIFO_blk[27] | proc_12_input_sync_blk[27] | proc_12_output_sync_blk[27]);
    assign proc_12_data_FIFO_blk[28] = 1'b0;
    assign proc_12_data_PIPO_blk[28] = 1'b0;
    assign proc_12_start_FIFO_blk[28] = 1'b0;
    assign proc_12_TLF_FIFO_blk[28] = 1'b0;
    assign proc_12_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_12_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_12[28] = dl_detect_out ? proc_dep_vld_vec_12_reg[28] : (proc_12_data_FIFO_blk[28] | proc_12_data_PIPO_blk[28] | proc_12_start_FIFO_blk[28] | proc_12_TLF_FIFO_blk[28] | proc_12_input_sync_blk[28] | proc_12_output_sync_blk[28]);
    assign proc_12_data_FIFO_blk[29] = 1'b0;
    assign proc_12_data_PIPO_blk[29] = 1'b0;
    assign proc_12_start_FIFO_blk[29] = 1'b0;
    assign proc_12_TLF_FIFO_blk[29] = 1'b0;
    assign proc_12_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_12_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_12[29] = dl_detect_out ? proc_dep_vld_vec_12_reg[29] : (proc_12_data_FIFO_blk[29] | proc_12_data_PIPO_blk[29] | proc_12_start_FIFO_blk[29] | proc_12_TLF_FIFO_blk[29] | proc_12_input_sync_blk[29] | proc_12_output_sync_blk[29]);
    assign proc_12_data_FIFO_blk[30] = 1'b0;
    assign proc_12_data_PIPO_blk[30] = 1'b0;
    assign proc_12_start_FIFO_blk[30] = 1'b0;
    assign proc_12_TLF_FIFO_blk[30] = 1'b0;
    assign proc_12_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_12_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_12[30] = dl_detect_out ? proc_dep_vld_vec_12_reg[30] : (proc_12_data_FIFO_blk[30] | proc_12_data_PIPO_blk[30] | proc_12_start_FIFO_blk[30] | proc_12_TLF_FIFO_blk[30] | proc_12_input_sync_blk[30] | proc_12_output_sync_blk[30]);
    assign proc_12_data_FIFO_blk[31] = 1'b0;
    assign proc_12_data_PIPO_blk[31] = 1'b0;
    assign proc_12_start_FIFO_blk[31] = 1'b0;
    assign proc_12_TLF_FIFO_blk[31] = 1'b0;
    assign proc_12_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_12_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_12[31] = dl_detect_out ? proc_dep_vld_vec_12_reg[31] : (proc_12_data_FIFO_blk[31] | proc_12_data_PIPO_blk[31] | proc_12_start_FIFO_blk[31] | proc_12_TLF_FIFO_blk[31] | proc_12_input_sync_blk[31] | proc_12_output_sync_blk[31]);
    assign proc_12_data_FIFO_blk[32] = 1'b0;
    assign proc_12_data_PIPO_blk[32] = 1'b0;
    assign proc_12_start_FIFO_blk[32] = 1'b0;
    assign proc_12_TLF_FIFO_blk[32] = 1'b0;
    assign proc_12_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_7_U0_ap_ready & ProcessingElement_7_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_12_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_12[32] = dl_detect_out ? proc_dep_vld_vec_12_reg[32] : (proc_12_data_FIFO_blk[32] | proc_12_data_PIPO_blk[32] | proc_12_start_FIFO_blk[32] | proc_12_TLF_FIFO_blk[32] | proc_12_input_sync_blk[32] | proc_12_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_12_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_12_reg <= proc_dep_vld_vec_12;
        end
    end
    assign in_chan_dep_vld_vec_12[0] = dep_chan_vld_0_12;
    assign in_chan_dep_data_vec_12[39 : 0] = dep_chan_data_0_12;
    assign token_in_vec_12[0] = token_0_12;
    assign in_chan_dep_vld_vec_12[1] = dep_chan_vld_1_12;
    assign in_chan_dep_data_vec_12[79 : 40] = dep_chan_data_1_12;
    assign token_in_vec_12[1] = token_1_12;
    assign in_chan_dep_vld_vec_12[2] = dep_chan_vld_3_12;
    assign in_chan_dep_data_vec_12[119 : 80] = dep_chan_data_3_12;
    assign token_in_vec_12[2] = token_3_12;
    assign in_chan_dep_vld_vec_12[3] = dep_chan_vld_6_12;
    assign in_chan_dep_data_vec_12[159 : 120] = dep_chan_data_6_12;
    assign token_in_vec_12[3] = token_6_12;
    assign in_chan_dep_vld_vec_12[4] = dep_chan_vld_7_12;
    assign in_chan_dep_data_vec_12[199 : 160] = dep_chan_data_7_12;
    assign token_in_vec_12[4] = token_7_12;
    assign in_chan_dep_vld_vec_12[5] = dep_chan_vld_8_12;
    assign in_chan_dep_data_vec_12[239 : 200] = dep_chan_data_8_12;
    assign token_in_vec_12[5] = token_8_12;
    assign in_chan_dep_vld_vec_12[6] = dep_chan_vld_9_12;
    assign in_chan_dep_data_vec_12[279 : 240] = dep_chan_data_9_12;
    assign token_in_vec_12[6] = token_9_12;
    assign in_chan_dep_vld_vec_12[7] = dep_chan_vld_10_12;
    assign in_chan_dep_data_vec_12[319 : 280] = dep_chan_data_10_12;
    assign token_in_vec_12[7] = token_10_12;
    assign in_chan_dep_vld_vec_12[8] = dep_chan_vld_11_12;
    assign in_chan_dep_data_vec_12[359 : 320] = dep_chan_data_11_12;
    assign token_in_vec_12[8] = token_11_12;
    assign in_chan_dep_vld_vec_12[9] = dep_chan_vld_13_12;
    assign in_chan_dep_data_vec_12[399 : 360] = dep_chan_data_13_12;
    assign token_in_vec_12[9] = token_13_12;
    assign in_chan_dep_vld_vec_12[10] = dep_chan_vld_14_12;
    assign in_chan_dep_data_vec_12[439 : 400] = dep_chan_data_14_12;
    assign token_in_vec_12[10] = token_14_12;
    assign in_chan_dep_vld_vec_12[11] = dep_chan_vld_15_12;
    assign in_chan_dep_data_vec_12[479 : 440] = dep_chan_data_15_12;
    assign token_in_vec_12[11] = token_15_12;
    assign in_chan_dep_vld_vec_12[12] = dep_chan_vld_16_12;
    assign in_chan_dep_data_vec_12[519 : 480] = dep_chan_data_16_12;
    assign token_in_vec_12[12] = token_16_12;
    assign in_chan_dep_vld_vec_12[13] = dep_chan_vld_17_12;
    assign in_chan_dep_data_vec_12[559 : 520] = dep_chan_data_17_12;
    assign token_in_vec_12[13] = token_17_12;
    assign in_chan_dep_vld_vec_12[14] = dep_chan_vld_18_12;
    assign in_chan_dep_data_vec_12[599 : 560] = dep_chan_data_18_12;
    assign token_in_vec_12[14] = token_18_12;
    assign in_chan_dep_vld_vec_12[15] = dep_chan_vld_19_12;
    assign in_chan_dep_data_vec_12[639 : 600] = dep_chan_data_19_12;
    assign token_in_vec_12[15] = token_19_12;
    assign in_chan_dep_vld_vec_12[16] = dep_chan_vld_20_12;
    assign in_chan_dep_data_vec_12[679 : 640] = dep_chan_data_20_12;
    assign token_in_vec_12[16] = token_20_12;
    assign in_chan_dep_vld_vec_12[17] = dep_chan_vld_21_12;
    assign in_chan_dep_data_vec_12[719 : 680] = dep_chan_data_21_12;
    assign token_in_vec_12[17] = token_21_12;
    assign in_chan_dep_vld_vec_12[18] = dep_chan_vld_22_12;
    assign in_chan_dep_data_vec_12[759 : 720] = dep_chan_data_22_12;
    assign token_in_vec_12[18] = token_22_12;
    assign in_chan_dep_vld_vec_12[19] = dep_chan_vld_23_12;
    assign in_chan_dep_data_vec_12[799 : 760] = dep_chan_data_23_12;
    assign token_in_vec_12[19] = token_23_12;
    assign in_chan_dep_vld_vec_12[20] = dep_chan_vld_24_12;
    assign in_chan_dep_data_vec_12[839 : 800] = dep_chan_data_24_12;
    assign token_in_vec_12[20] = token_24_12;
    assign in_chan_dep_vld_vec_12[21] = dep_chan_vld_25_12;
    assign in_chan_dep_data_vec_12[879 : 840] = dep_chan_data_25_12;
    assign token_in_vec_12[21] = token_25_12;
    assign in_chan_dep_vld_vec_12[22] = dep_chan_vld_26_12;
    assign in_chan_dep_data_vec_12[919 : 880] = dep_chan_data_26_12;
    assign token_in_vec_12[22] = token_26_12;
    assign in_chan_dep_vld_vec_12[23] = dep_chan_vld_27_12;
    assign in_chan_dep_data_vec_12[959 : 920] = dep_chan_data_27_12;
    assign token_in_vec_12[23] = token_27_12;
    assign in_chan_dep_vld_vec_12[24] = dep_chan_vld_28_12;
    assign in_chan_dep_data_vec_12[999 : 960] = dep_chan_data_28_12;
    assign token_in_vec_12[24] = token_28_12;
    assign in_chan_dep_vld_vec_12[25] = dep_chan_vld_29_12;
    assign in_chan_dep_data_vec_12[1039 : 1000] = dep_chan_data_29_12;
    assign token_in_vec_12[25] = token_29_12;
    assign in_chan_dep_vld_vec_12[26] = dep_chan_vld_30_12;
    assign in_chan_dep_data_vec_12[1079 : 1040] = dep_chan_data_30_12;
    assign token_in_vec_12[26] = token_30_12;
    assign in_chan_dep_vld_vec_12[27] = dep_chan_vld_31_12;
    assign in_chan_dep_data_vec_12[1119 : 1080] = dep_chan_data_31_12;
    assign token_in_vec_12[27] = token_31_12;
    assign in_chan_dep_vld_vec_12[28] = dep_chan_vld_32_12;
    assign in_chan_dep_data_vec_12[1159 : 1120] = dep_chan_data_32_12;
    assign token_in_vec_12[28] = token_32_12;
    assign in_chan_dep_vld_vec_12[29] = dep_chan_vld_33_12;
    assign in_chan_dep_data_vec_12[1199 : 1160] = dep_chan_data_33_12;
    assign token_in_vec_12[29] = token_33_12;
    assign in_chan_dep_vld_vec_12[30] = dep_chan_vld_34_12;
    assign in_chan_dep_data_vec_12[1239 : 1200] = dep_chan_data_34_12;
    assign token_in_vec_12[30] = token_34_12;
    assign in_chan_dep_vld_vec_12[31] = dep_chan_vld_35_12;
    assign in_chan_dep_data_vec_12[1279 : 1240] = dep_chan_data_35_12;
    assign token_in_vec_12[31] = token_35_12;
    assign in_chan_dep_vld_vec_12[32] = dep_chan_vld_36_12;
    assign in_chan_dep_data_vec_12[1319 : 1280] = dep_chan_data_36_12;
    assign token_in_vec_12[32] = token_36_12;
    assign dep_chan_vld_12_11 = out_chan_dep_vld_vec_12[0];
    assign dep_chan_data_12_11 = out_chan_dep_data_12;
    assign token_12_11 = token_out_vec_12[0];
    assign dep_chan_vld_12_13 = out_chan_dep_vld_vec_12[1];
    assign dep_chan_data_12_13 = out_chan_dep_data_12;
    assign token_12_13 = token_out_vec_12[1];
    assign dep_chan_vld_12_0 = out_chan_dep_vld_vec_12[2];
    assign dep_chan_data_12_0 = out_chan_dep_data_12;
    assign token_12_0 = token_out_vec_12[2];
    assign dep_chan_vld_12_1 = out_chan_dep_vld_vec_12[3];
    assign dep_chan_data_12_1 = out_chan_dep_data_12;
    assign token_12_1 = token_out_vec_12[3];
    assign dep_chan_vld_12_3 = out_chan_dep_vld_vec_12[4];
    assign dep_chan_data_12_3 = out_chan_dep_data_12;
    assign token_12_3 = token_out_vec_12[4];
    assign dep_chan_vld_12_6 = out_chan_dep_vld_vec_12[5];
    assign dep_chan_data_12_6 = out_chan_dep_data_12;
    assign token_12_6 = token_out_vec_12[5];
    assign dep_chan_vld_12_7 = out_chan_dep_vld_vec_12[6];
    assign dep_chan_data_12_7 = out_chan_dep_data_12;
    assign token_12_7 = token_out_vec_12[6];
    assign dep_chan_vld_12_8 = out_chan_dep_vld_vec_12[7];
    assign dep_chan_data_12_8 = out_chan_dep_data_12;
    assign token_12_8 = token_out_vec_12[7];
    assign dep_chan_vld_12_9 = out_chan_dep_vld_vec_12[8];
    assign dep_chan_data_12_9 = out_chan_dep_data_12;
    assign token_12_9 = token_out_vec_12[8];
    assign dep_chan_vld_12_10 = out_chan_dep_vld_vec_12[9];
    assign dep_chan_data_12_10 = out_chan_dep_data_12;
    assign token_12_10 = token_out_vec_12[9];
    assign dep_chan_vld_12_14 = out_chan_dep_vld_vec_12[10];
    assign dep_chan_data_12_14 = out_chan_dep_data_12;
    assign token_12_14 = token_out_vec_12[10];
    assign dep_chan_vld_12_15 = out_chan_dep_vld_vec_12[11];
    assign dep_chan_data_12_15 = out_chan_dep_data_12;
    assign token_12_15 = token_out_vec_12[11];
    assign dep_chan_vld_12_16 = out_chan_dep_vld_vec_12[12];
    assign dep_chan_data_12_16 = out_chan_dep_data_12;
    assign token_12_16 = token_out_vec_12[12];
    assign dep_chan_vld_12_17 = out_chan_dep_vld_vec_12[13];
    assign dep_chan_data_12_17 = out_chan_dep_data_12;
    assign token_12_17 = token_out_vec_12[13];
    assign dep_chan_vld_12_18 = out_chan_dep_vld_vec_12[14];
    assign dep_chan_data_12_18 = out_chan_dep_data_12;
    assign token_12_18 = token_out_vec_12[14];
    assign dep_chan_vld_12_19 = out_chan_dep_vld_vec_12[15];
    assign dep_chan_data_12_19 = out_chan_dep_data_12;
    assign token_12_19 = token_out_vec_12[15];
    assign dep_chan_vld_12_20 = out_chan_dep_vld_vec_12[16];
    assign dep_chan_data_12_20 = out_chan_dep_data_12;
    assign token_12_20 = token_out_vec_12[16];
    assign dep_chan_vld_12_21 = out_chan_dep_vld_vec_12[17];
    assign dep_chan_data_12_21 = out_chan_dep_data_12;
    assign token_12_21 = token_out_vec_12[17];
    assign dep_chan_vld_12_22 = out_chan_dep_vld_vec_12[18];
    assign dep_chan_data_12_22 = out_chan_dep_data_12;
    assign token_12_22 = token_out_vec_12[18];
    assign dep_chan_vld_12_23 = out_chan_dep_vld_vec_12[19];
    assign dep_chan_data_12_23 = out_chan_dep_data_12;
    assign token_12_23 = token_out_vec_12[19];
    assign dep_chan_vld_12_24 = out_chan_dep_vld_vec_12[20];
    assign dep_chan_data_12_24 = out_chan_dep_data_12;
    assign token_12_24 = token_out_vec_12[20];
    assign dep_chan_vld_12_25 = out_chan_dep_vld_vec_12[21];
    assign dep_chan_data_12_25 = out_chan_dep_data_12;
    assign token_12_25 = token_out_vec_12[21];
    assign dep_chan_vld_12_26 = out_chan_dep_vld_vec_12[22];
    assign dep_chan_data_12_26 = out_chan_dep_data_12;
    assign token_12_26 = token_out_vec_12[22];
    assign dep_chan_vld_12_27 = out_chan_dep_vld_vec_12[23];
    assign dep_chan_data_12_27 = out_chan_dep_data_12;
    assign token_12_27 = token_out_vec_12[23];
    assign dep_chan_vld_12_28 = out_chan_dep_vld_vec_12[24];
    assign dep_chan_data_12_28 = out_chan_dep_data_12;
    assign token_12_28 = token_out_vec_12[24];
    assign dep_chan_vld_12_29 = out_chan_dep_vld_vec_12[25];
    assign dep_chan_data_12_29 = out_chan_dep_data_12;
    assign token_12_29 = token_out_vec_12[25];
    assign dep_chan_vld_12_30 = out_chan_dep_vld_vec_12[26];
    assign dep_chan_data_12_30 = out_chan_dep_data_12;
    assign token_12_30 = token_out_vec_12[26];
    assign dep_chan_vld_12_31 = out_chan_dep_vld_vec_12[27];
    assign dep_chan_data_12_31 = out_chan_dep_data_12;
    assign token_12_31 = token_out_vec_12[27];
    assign dep_chan_vld_12_32 = out_chan_dep_vld_vec_12[28];
    assign dep_chan_data_12_32 = out_chan_dep_data_12;
    assign token_12_32 = token_out_vec_12[28];
    assign dep_chan_vld_12_33 = out_chan_dep_vld_vec_12[29];
    assign dep_chan_data_12_33 = out_chan_dep_data_12;
    assign token_12_33 = token_out_vec_12[29];
    assign dep_chan_vld_12_34 = out_chan_dep_vld_vec_12[30];
    assign dep_chan_data_12_34 = out_chan_dep_data_12;
    assign token_12_34 = token_out_vec_12[30];
    assign dep_chan_vld_12_35 = out_chan_dep_vld_vec_12[31];
    assign dep_chan_data_12_35 = out_chan_dep_data_12;
    assign token_12_35 = token_out_vec_12[31];
    assign dep_chan_vld_12_36 = out_chan_dep_vld_vec_12[32];
    assign dep_chan_data_12_36 = out_chan_dep_data_12;
    assign token_12_36 = token_out_vec_12[32];

    // Process: ProcessingElement_8_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 13, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_13 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_13),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_13),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_13),
        .token_in_vec(token_in_vec_13),
        .dl_detect_in(dl_detect_out),
        .origin(origin[13]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_13),
        .out_chan_dep_data(out_chan_dep_data_13),
        .token_out_vec(token_out_vec_13),
        .dl_detect_out(dl_in_vec[13]));

    assign proc_13_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_7_blk_n) | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_7_blk_n) | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_WriteC_Flattened_fu_179.cPipes_7_blk_n);
    assign proc_13_data_PIPO_blk[0] = 1'b0;
    assign proc_13_start_FIFO_blk[0] = 1'b0;
    assign proc_13_TLF_FIFO_blk[0] = 1'b0;
    assign proc_13_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_13_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_13[0] = dl_detect_out ? proc_dep_vld_vec_13_reg[0] : (proc_13_data_FIFO_blk[0] | proc_13_data_PIPO_blk[0] | proc_13_start_FIFO_blk[0] | proc_13_TLF_FIFO_blk[0] | proc_13_input_sync_blk[0] | proc_13_output_sync_blk[0]);
    assign proc_13_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_8_blk_n) | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_8_blk_n) | (~ProcessingElement_8_U0.grp_ProcessingElement_8_Pipeline_WriteC_Flattened_fu_179.cPipes_8_blk_n);
    assign proc_13_data_PIPO_blk[1] = 1'b0;
    assign proc_13_start_FIFO_blk[1] = 1'b0;
    assign proc_13_TLF_FIFO_blk[1] = 1'b0;
    assign proc_13_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_13_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_13[1] = dl_detect_out ? proc_dep_vld_vec_13_reg[1] : (proc_13_data_FIFO_blk[1] | proc_13_data_PIPO_blk[1] | proc_13_start_FIFO_blk[1] | proc_13_TLF_FIFO_blk[1] | proc_13_input_sync_blk[1] | proc_13_output_sync_blk[1]);
    assign proc_13_data_FIFO_blk[2] = 1'b0;
    assign proc_13_data_PIPO_blk[2] = 1'b0;
    assign proc_13_start_FIFO_blk[2] = 1'b0;
    assign proc_13_TLF_FIFO_blk[2] = 1'b0;
    assign proc_13_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_13_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_13[2] = dl_detect_out ? proc_dep_vld_vec_13_reg[2] : (proc_13_data_FIFO_blk[2] | proc_13_data_PIPO_blk[2] | proc_13_start_FIFO_blk[2] | proc_13_TLF_FIFO_blk[2] | proc_13_input_sync_blk[2] | proc_13_output_sync_blk[2]);
    assign proc_13_data_FIFO_blk[3] = 1'b0;
    assign proc_13_data_PIPO_blk[3] = 1'b0;
    assign proc_13_start_FIFO_blk[3] = 1'b0;
    assign proc_13_TLF_FIFO_blk[3] = 1'b0;
    assign proc_13_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_13_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_13[3] = dl_detect_out ? proc_dep_vld_vec_13_reg[3] : (proc_13_data_FIFO_blk[3] | proc_13_data_PIPO_blk[3] | proc_13_start_FIFO_blk[3] | proc_13_TLF_FIFO_blk[3] | proc_13_input_sync_blk[3] | proc_13_output_sync_blk[3]);
    assign proc_13_data_FIFO_blk[4] = 1'b0;
    assign proc_13_data_PIPO_blk[4] = 1'b0;
    assign proc_13_start_FIFO_blk[4] = 1'b0;
    assign proc_13_TLF_FIFO_blk[4] = 1'b0;
    assign proc_13_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_13_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_13[4] = dl_detect_out ? proc_dep_vld_vec_13_reg[4] : (proc_13_data_FIFO_blk[4] | proc_13_data_PIPO_blk[4] | proc_13_start_FIFO_blk[4] | proc_13_TLF_FIFO_blk[4] | proc_13_input_sync_blk[4] | proc_13_output_sync_blk[4]);
    assign proc_13_data_FIFO_blk[5] = 1'b0;
    assign proc_13_data_PIPO_blk[5] = 1'b0;
    assign proc_13_start_FIFO_blk[5] = 1'b0;
    assign proc_13_TLF_FIFO_blk[5] = 1'b0;
    assign proc_13_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_13_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_13[5] = dl_detect_out ? proc_dep_vld_vec_13_reg[5] : (proc_13_data_FIFO_blk[5] | proc_13_data_PIPO_blk[5] | proc_13_start_FIFO_blk[5] | proc_13_TLF_FIFO_blk[5] | proc_13_input_sync_blk[5] | proc_13_output_sync_blk[5]);
    assign proc_13_data_FIFO_blk[6] = 1'b0;
    assign proc_13_data_PIPO_blk[6] = 1'b0;
    assign proc_13_start_FIFO_blk[6] = 1'b0;
    assign proc_13_TLF_FIFO_blk[6] = 1'b0;
    assign proc_13_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_13_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_13[6] = dl_detect_out ? proc_dep_vld_vec_13_reg[6] : (proc_13_data_FIFO_blk[6] | proc_13_data_PIPO_blk[6] | proc_13_start_FIFO_blk[6] | proc_13_TLF_FIFO_blk[6] | proc_13_input_sync_blk[6] | proc_13_output_sync_blk[6]);
    assign proc_13_data_FIFO_blk[7] = 1'b0;
    assign proc_13_data_PIPO_blk[7] = 1'b0;
    assign proc_13_start_FIFO_blk[7] = 1'b0;
    assign proc_13_TLF_FIFO_blk[7] = 1'b0;
    assign proc_13_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_13_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_13[7] = dl_detect_out ? proc_dep_vld_vec_13_reg[7] : (proc_13_data_FIFO_blk[7] | proc_13_data_PIPO_blk[7] | proc_13_start_FIFO_blk[7] | proc_13_TLF_FIFO_blk[7] | proc_13_input_sync_blk[7] | proc_13_output_sync_blk[7]);
    assign proc_13_data_FIFO_blk[8] = 1'b0;
    assign proc_13_data_PIPO_blk[8] = 1'b0;
    assign proc_13_start_FIFO_blk[8] = 1'b0;
    assign proc_13_TLF_FIFO_blk[8] = 1'b0;
    assign proc_13_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_13_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_13[8] = dl_detect_out ? proc_dep_vld_vec_13_reg[8] : (proc_13_data_FIFO_blk[8] | proc_13_data_PIPO_blk[8] | proc_13_start_FIFO_blk[8] | proc_13_TLF_FIFO_blk[8] | proc_13_input_sync_blk[8] | proc_13_output_sync_blk[8]);
    assign proc_13_data_FIFO_blk[9] = 1'b0;
    assign proc_13_data_PIPO_blk[9] = 1'b0;
    assign proc_13_start_FIFO_blk[9] = 1'b0;
    assign proc_13_TLF_FIFO_blk[9] = 1'b0;
    assign proc_13_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_13_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_13[9] = dl_detect_out ? proc_dep_vld_vec_13_reg[9] : (proc_13_data_FIFO_blk[9] | proc_13_data_PIPO_blk[9] | proc_13_start_FIFO_blk[9] | proc_13_TLF_FIFO_blk[9] | proc_13_input_sync_blk[9] | proc_13_output_sync_blk[9]);
    assign proc_13_data_FIFO_blk[10] = 1'b0;
    assign proc_13_data_PIPO_blk[10] = 1'b0;
    assign proc_13_start_FIFO_blk[10] = 1'b0;
    assign proc_13_TLF_FIFO_blk[10] = 1'b0;
    assign proc_13_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_13_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_13[10] = dl_detect_out ? proc_dep_vld_vec_13_reg[10] : (proc_13_data_FIFO_blk[10] | proc_13_data_PIPO_blk[10] | proc_13_start_FIFO_blk[10] | proc_13_TLF_FIFO_blk[10] | proc_13_input_sync_blk[10] | proc_13_output_sync_blk[10]);
    assign proc_13_data_FIFO_blk[11] = 1'b0;
    assign proc_13_data_PIPO_blk[11] = 1'b0;
    assign proc_13_start_FIFO_blk[11] = 1'b0;
    assign proc_13_TLF_FIFO_blk[11] = 1'b0;
    assign proc_13_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_13_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_13[11] = dl_detect_out ? proc_dep_vld_vec_13_reg[11] : (proc_13_data_FIFO_blk[11] | proc_13_data_PIPO_blk[11] | proc_13_start_FIFO_blk[11] | proc_13_TLF_FIFO_blk[11] | proc_13_input_sync_blk[11] | proc_13_output_sync_blk[11]);
    assign proc_13_data_FIFO_blk[12] = 1'b0;
    assign proc_13_data_PIPO_blk[12] = 1'b0;
    assign proc_13_start_FIFO_blk[12] = 1'b0;
    assign proc_13_TLF_FIFO_blk[12] = 1'b0;
    assign proc_13_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_13_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_13[12] = dl_detect_out ? proc_dep_vld_vec_13_reg[12] : (proc_13_data_FIFO_blk[12] | proc_13_data_PIPO_blk[12] | proc_13_start_FIFO_blk[12] | proc_13_TLF_FIFO_blk[12] | proc_13_input_sync_blk[12] | proc_13_output_sync_blk[12]);
    assign proc_13_data_FIFO_blk[13] = 1'b0;
    assign proc_13_data_PIPO_blk[13] = 1'b0;
    assign proc_13_start_FIFO_blk[13] = 1'b0;
    assign proc_13_TLF_FIFO_blk[13] = 1'b0;
    assign proc_13_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_13_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_13[13] = dl_detect_out ? proc_dep_vld_vec_13_reg[13] : (proc_13_data_FIFO_blk[13] | proc_13_data_PIPO_blk[13] | proc_13_start_FIFO_blk[13] | proc_13_TLF_FIFO_blk[13] | proc_13_input_sync_blk[13] | proc_13_output_sync_blk[13]);
    assign proc_13_data_FIFO_blk[14] = 1'b0;
    assign proc_13_data_PIPO_blk[14] = 1'b0;
    assign proc_13_start_FIFO_blk[14] = 1'b0;
    assign proc_13_TLF_FIFO_blk[14] = 1'b0;
    assign proc_13_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_13_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_13[14] = dl_detect_out ? proc_dep_vld_vec_13_reg[14] : (proc_13_data_FIFO_blk[14] | proc_13_data_PIPO_blk[14] | proc_13_start_FIFO_blk[14] | proc_13_TLF_FIFO_blk[14] | proc_13_input_sync_blk[14] | proc_13_output_sync_blk[14]);
    assign proc_13_data_FIFO_blk[15] = 1'b0;
    assign proc_13_data_PIPO_blk[15] = 1'b0;
    assign proc_13_start_FIFO_blk[15] = 1'b0;
    assign proc_13_TLF_FIFO_blk[15] = 1'b0;
    assign proc_13_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_13_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_13[15] = dl_detect_out ? proc_dep_vld_vec_13_reg[15] : (proc_13_data_FIFO_blk[15] | proc_13_data_PIPO_blk[15] | proc_13_start_FIFO_blk[15] | proc_13_TLF_FIFO_blk[15] | proc_13_input_sync_blk[15] | proc_13_output_sync_blk[15]);
    assign proc_13_data_FIFO_blk[16] = 1'b0;
    assign proc_13_data_PIPO_blk[16] = 1'b0;
    assign proc_13_start_FIFO_blk[16] = 1'b0;
    assign proc_13_TLF_FIFO_blk[16] = 1'b0;
    assign proc_13_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_13_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_13[16] = dl_detect_out ? proc_dep_vld_vec_13_reg[16] : (proc_13_data_FIFO_blk[16] | proc_13_data_PIPO_blk[16] | proc_13_start_FIFO_blk[16] | proc_13_TLF_FIFO_blk[16] | proc_13_input_sync_blk[16] | proc_13_output_sync_blk[16]);
    assign proc_13_data_FIFO_blk[17] = 1'b0;
    assign proc_13_data_PIPO_blk[17] = 1'b0;
    assign proc_13_start_FIFO_blk[17] = 1'b0;
    assign proc_13_TLF_FIFO_blk[17] = 1'b0;
    assign proc_13_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_13_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_13[17] = dl_detect_out ? proc_dep_vld_vec_13_reg[17] : (proc_13_data_FIFO_blk[17] | proc_13_data_PIPO_blk[17] | proc_13_start_FIFO_blk[17] | proc_13_TLF_FIFO_blk[17] | proc_13_input_sync_blk[17] | proc_13_output_sync_blk[17]);
    assign proc_13_data_FIFO_blk[18] = 1'b0;
    assign proc_13_data_PIPO_blk[18] = 1'b0;
    assign proc_13_start_FIFO_blk[18] = 1'b0;
    assign proc_13_TLF_FIFO_blk[18] = 1'b0;
    assign proc_13_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_13_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_13[18] = dl_detect_out ? proc_dep_vld_vec_13_reg[18] : (proc_13_data_FIFO_blk[18] | proc_13_data_PIPO_blk[18] | proc_13_start_FIFO_blk[18] | proc_13_TLF_FIFO_blk[18] | proc_13_input_sync_blk[18] | proc_13_output_sync_blk[18]);
    assign proc_13_data_FIFO_blk[19] = 1'b0;
    assign proc_13_data_PIPO_blk[19] = 1'b0;
    assign proc_13_start_FIFO_blk[19] = 1'b0;
    assign proc_13_TLF_FIFO_blk[19] = 1'b0;
    assign proc_13_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_13_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_13[19] = dl_detect_out ? proc_dep_vld_vec_13_reg[19] : (proc_13_data_FIFO_blk[19] | proc_13_data_PIPO_blk[19] | proc_13_start_FIFO_blk[19] | proc_13_TLF_FIFO_blk[19] | proc_13_input_sync_blk[19] | proc_13_output_sync_blk[19]);
    assign proc_13_data_FIFO_blk[20] = 1'b0;
    assign proc_13_data_PIPO_blk[20] = 1'b0;
    assign proc_13_start_FIFO_blk[20] = 1'b0;
    assign proc_13_TLF_FIFO_blk[20] = 1'b0;
    assign proc_13_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_13_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_13[20] = dl_detect_out ? proc_dep_vld_vec_13_reg[20] : (proc_13_data_FIFO_blk[20] | proc_13_data_PIPO_blk[20] | proc_13_start_FIFO_blk[20] | proc_13_TLF_FIFO_blk[20] | proc_13_input_sync_blk[20] | proc_13_output_sync_blk[20]);
    assign proc_13_data_FIFO_blk[21] = 1'b0;
    assign proc_13_data_PIPO_blk[21] = 1'b0;
    assign proc_13_start_FIFO_blk[21] = 1'b0;
    assign proc_13_TLF_FIFO_blk[21] = 1'b0;
    assign proc_13_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_13_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_13[21] = dl_detect_out ? proc_dep_vld_vec_13_reg[21] : (proc_13_data_FIFO_blk[21] | proc_13_data_PIPO_blk[21] | proc_13_start_FIFO_blk[21] | proc_13_TLF_FIFO_blk[21] | proc_13_input_sync_blk[21] | proc_13_output_sync_blk[21]);
    assign proc_13_data_FIFO_blk[22] = 1'b0;
    assign proc_13_data_PIPO_blk[22] = 1'b0;
    assign proc_13_start_FIFO_blk[22] = 1'b0;
    assign proc_13_TLF_FIFO_blk[22] = 1'b0;
    assign proc_13_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_13_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_13[22] = dl_detect_out ? proc_dep_vld_vec_13_reg[22] : (proc_13_data_FIFO_blk[22] | proc_13_data_PIPO_blk[22] | proc_13_start_FIFO_blk[22] | proc_13_TLF_FIFO_blk[22] | proc_13_input_sync_blk[22] | proc_13_output_sync_blk[22]);
    assign proc_13_data_FIFO_blk[23] = 1'b0;
    assign proc_13_data_PIPO_blk[23] = 1'b0;
    assign proc_13_start_FIFO_blk[23] = 1'b0;
    assign proc_13_TLF_FIFO_blk[23] = 1'b0;
    assign proc_13_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_13_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_13[23] = dl_detect_out ? proc_dep_vld_vec_13_reg[23] : (proc_13_data_FIFO_blk[23] | proc_13_data_PIPO_blk[23] | proc_13_start_FIFO_blk[23] | proc_13_TLF_FIFO_blk[23] | proc_13_input_sync_blk[23] | proc_13_output_sync_blk[23]);
    assign proc_13_data_FIFO_blk[24] = 1'b0;
    assign proc_13_data_PIPO_blk[24] = 1'b0;
    assign proc_13_start_FIFO_blk[24] = 1'b0;
    assign proc_13_TLF_FIFO_blk[24] = 1'b0;
    assign proc_13_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_13_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_13[24] = dl_detect_out ? proc_dep_vld_vec_13_reg[24] : (proc_13_data_FIFO_blk[24] | proc_13_data_PIPO_blk[24] | proc_13_start_FIFO_blk[24] | proc_13_TLF_FIFO_blk[24] | proc_13_input_sync_blk[24] | proc_13_output_sync_blk[24]);
    assign proc_13_data_FIFO_blk[25] = 1'b0;
    assign proc_13_data_PIPO_blk[25] = 1'b0;
    assign proc_13_start_FIFO_blk[25] = 1'b0;
    assign proc_13_TLF_FIFO_blk[25] = 1'b0;
    assign proc_13_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_13_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_13[25] = dl_detect_out ? proc_dep_vld_vec_13_reg[25] : (proc_13_data_FIFO_blk[25] | proc_13_data_PIPO_blk[25] | proc_13_start_FIFO_blk[25] | proc_13_TLF_FIFO_blk[25] | proc_13_input_sync_blk[25] | proc_13_output_sync_blk[25]);
    assign proc_13_data_FIFO_blk[26] = 1'b0;
    assign proc_13_data_PIPO_blk[26] = 1'b0;
    assign proc_13_start_FIFO_blk[26] = 1'b0;
    assign proc_13_TLF_FIFO_blk[26] = 1'b0;
    assign proc_13_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_13_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_13[26] = dl_detect_out ? proc_dep_vld_vec_13_reg[26] : (proc_13_data_FIFO_blk[26] | proc_13_data_PIPO_blk[26] | proc_13_start_FIFO_blk[26] | proc_13_TLF_FIFO_blk[26] | proc_13_input_sync_blk[26] | proc_13_output_sync_blk[26]);
    assign proc_13_data_FIFO_blk[27] = 1'b0;
    assign proc_13_data_PIPO_blk[27] = 1'b0;
    assign proc_13_start_FIFO_blk[27] = 1'b0;
    assign proc_13_TLF_FIFO_blk[27] = 1'b0;
    assign proc_13_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_13_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_13[27] = dl_detect_out ? proc_dep_vld_vec_13_reg[27] : (proc_13_data_FIFO_blk[27] | proc_13_data_PIPO_blk[27] | proc_13_start_FIFO_blk[27] | proc_13_TLF_FIFO_blk[27] | proc_13_input_sync_blk[27] | proc_13_output_sync_blk[27]);
    assign proc_13_data_FIFO_blk[28] = 1'b0;
    assign proc_13_data_PIPO_blk[28] = 1'b0;
    assign proc_13_start_FIFO_blk[28] = 1'b0;
    assign proc_13_TLF_FIFO_blk[28] = 1'b0;
    assign proc_13_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_13_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_13[28] = dl_detect_out ? proc_dep_vld_vec_13_reg[28] : (proc_13_data_FIFO_blk[28] | proc_13_data_PIPO_blk[28] | proc_13_start_FIFO_blk[28] | proc_13_TLF_FIFO_blk[28] | proc_13_input_sync_blk[28] | proc_13_output_sync_blk[28]);
    assign proc_13_data_FIFO_blk[29] = 1'b0;
    assign proc_13_data_PIPO_blk[29] = 1'b0;
    assign proc_13_start_FIFO_blk[29] = 1'b0;
    assign proc_13_TLF_FIFO_blk[29] = 1'b0;
    assign proc_13_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_13_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_13[29] = dl_detect_out ? proc_dep_vld_vec_13_reg[29] : (proc_13_data_FIFO_blk[29] | proc_13_data_PIPO_blk[29] | proc_13_start_FIFO_blk[29] | proc_13_TLF_FIFO_blk[29] | proc_13_input_sync_blk[29] | proc_13_output_sync_blk[29]);
    assign proc_13_data_FIFO_blk[30] = 1'b0;
    assign proc_13_data_PIPO_blk[30] = 1'b0;
    assign proc_13_start_FIFO_blk[30] = 1'b0;
    assign proc_13_TLF_FIFO_blk[30] = 1'b0;
    assign proc_13_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_13_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_13[30] = dl_detect_out ? proc_dep_vld_vec_13_reg[30] : (proc_13_data_FIFO_blk[30] | proc_13_data_PIPO_blk[30] | proc_13_start_FIFO_blk[30] | proc_13_TLF_FIFO_blk[30] | proc_13_input_sync_blk[30] | proc_13_output_sync_blk[30]);
    assign proc_13_data_FIFO_blk[31] = 1'b0;
    assign proc_13_data_PIPO_blk[31] = 1'b0;
    assign proc_13_start_FIFO_blk[31] = 1'b0;
    assign proc_13_TLF_FIFO_blk[31] = 1'b0;
    assign proc_13_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_13_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_13[31] = dl_detect_out ? proc_dep_vld_vec_13_reg[31] : (proc_13_data_FIFO_blk[31] | proc_13_data_PIPO_blk[31] | proc_13_start_FIFO_blk[31] | proc_13_TLF_FIFO_blk[31] | proc_13_input_sync_blk[31] | proc_13_output_sync_blk[31]);
    assign proc_13_data_FIFO_blk[32] = 1'b0;
    assign proc_13_data_PIPO_blk[32] = 1'b0;
    assign proc_13_start_FIFO_blk[32] = 1'b0;
    assign proc_13_TLF_FIFO_blk[32] = 1'b0;
    assign proc_13_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_8_U0_ap_ready & ProcessingElement_8_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_13_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_13[32] = dl_detect_out ? proc_dep_vld_vec_13_reg[32] : (proc_13_data_FIFO_blk[32] | proc_13_data_PIPO_blk[32] | proc_13_start_FIFO_blk[32] | proc_13_TLF_FIFO_blk[32] | proc_13_input_sync_blk[32] | proc_13_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_13_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_13_reg <= proc_dep_vld_vec_13;
        end
    end
    assign in_chan_dep_vld_vec_13[0] = dep_chan_vld_0_13;
    assign in_chan_dep_data_vec_13[39 : 0] = dep_chan_data_0_13;
    assign token_in_vec_13[0] = token_0_13;
    assign in_chan_dep_vld_vec_13[1] = dep_chan_vld_1_13;
    assign in_chan_dep_data_vec_13[79 : 40] = dep_chan_data_1_13;
    assign token_in_vec_13[1] = token_1_13;
    assign in_chan_dep_vld_vec_13[2] = dep_chan_vld_3_13;
    assign in_chan_dep_data_vec_13[119 : 80] = dep_chan_data_3_13;
    assign token_in_vec_13[2] = token_3_13;
    assign in_chan_dep_vld_vec_13[3] = dep_chan_vld_6_13;
    assign in_chan_dep_data_vec_13[159 : 120] = dep_chan_data_6_13;
    assign token_in_vec_13[3] = token_6_13;
    assign in_chan_dep_vld_vec_13[4] = dep_chan_vld_7_13;
    assign in_chan_dep_data_vec_13[199 : 160] = dep_chan_data_7_13;
    assign token_in_vec_13[4] = token_7_13;
    assign in_chan_dep_vld_vec_13[5] = dep_chan_vld_8_13;
    assign in_chan_dep_data_vec_13[239 : 200] = dep_chan_data_8_13;
    assign token_in_vec_13[5] = token_8_13;
    assign in_chan_dep_vld_vec_13[6] = dep_chan_vld_9_13;
    assign in_chan_dep_data_vec_13[279 : 240] = dep_chan_data_9_13;
    assign token_in_vec_13[6] = token_9_13;
    assign in_chan_dep_vld_vec_13[7] = dep_chan_vld_10_13;
    assign in_chan_dep_data_vec_13[319 : 280] = dep_chan_data_10_13;
    assign token_in_vec_13[7] = token_10_13;
    assign in_chan_dep_vld_vec_13[8] = dep_chan_vld_11_13;
    assign in_chan_dep_data_vec_13[359 : 320] = dep_chan_data_11_13;
    assign token_in_vec_13[8] = token_11_13;
    assign in_chan_dep_vld_vec_13[9] = dep_chan_vld_12_13;
    assign in_chan_dep_data_vec_13[399 : 360] = dep_chan_data_12_13;
    assign token_in_vec_13[9] = token_12_13;
    assign in_chan_dep_vld_vec_13[10] = dep_chan_vld_14_13;
    assign in_chan_dep_data_vec_13[439 : 400] = dep_chan_data_14_13;
    assign token_in_vec_13[10] = token_14_13;
    assign in_chan_dep_vld_vec_13[11] = dep_chan_vld_15_13;
    assign in_chan_dep_data_vec_13[479 : 440] = dep_chan_data_15_13;
    assign token_in_vec_13[11] = token_15_13;
    assign in_chan_dep_vld_vec_13[12] = dep_chan_vld_16_13;
    assign in_chan_dep_data_vec_13[519 : 480] = dep_chan_data_16_13;
    assign token_in_vec_13[12] = token_16_13;
    assign in_chan_dep_vld_vec_13[13] = dep_chan_vld_17_13;
    assign in_chan_dep_data_vec_13[559 : 520] = dep_chan_data_17_13;
    assign token_in_vec_13[13] = token_17_13;
    assign in_chan_dep_vld_vec_13[14] = dep_chan_vld_18_13;
    assign in_chan_dep_data_vec_13[599 : 560] = dep_chan_data_18_13;
    assign token_in_vec_13[14] = token_18_13;
    assign in_chan_dep_vld_vec_13[15] = dep_chan_vld_19_13;
    assign in_chan_dep_data_vec_13[639 : 600] = dep_chan_data_19_13;
    assign token_in_vec_13[15] = token_19_13;
    assign in_chan_dep_vld_vec_13[16] = dep_chan_vld_20_13;
    assign in_chan_dep_data_vec_13[679 : 640] = dep_chan_data_20_13;
    assign token_in_vec_13[16] = token_20_13;
    assign in_chan_dep_vld_vec_13[17] = dep_chan_vld_21_13;
    assign in_chan_dep_data_vec_13[719 : 680] = dep_chan_data_21_13;
    assign token_in_vec_13[17] = token_21_13;
    assign in_chan_dep_vld_vec_13[18] = dep_chan_vld_22_13;
    assign in_chan_dep_data_vec_13[759 : 720] = dep_chan_data_22_13;
    assign token_in_vec_13[18] = token_22_13;
    assign in_chan_dep_vld_vec_13[19] = dep_chan_vld_23_13;
    assign in_chan_dep_data_vec_13[799 : 760] = dep_chan_data_23_13;
    assign token_in_vec_13[19] = token_23_13;
    assign in_chan_dep_vld_vec_13[20] = dep_chan_vld_24_13;
    assign in_chan_dep_data_vec_13[839 : 800] = dep_chan_data_24_13;
    assign token_in_vec_13[20] = token_24_13;
    assign in_chan_dep_vld_vec_13[21] = dep_chan_vld_25_13;
    assign in_chan_dep_data_vec_13[879 : 840] = dep_chan_data_25_13;
    assign token_in_vec_13[21] = token_25_13;
    assign in_chan_dep_vld_vec_13[22] = dep_chan_vld_26_13;
    assign in_chan_dep_data_vec_13[919 : 880] = dep_chan_data_26_13;
    assign token_in_vec_13[22] = token_26_13;
    assign in_chan_dep_vld_vec_13[23] = dep_chan_vld_27_13;
    assign in_chan_dep_data_vec_13[959 : 920] = dep_chan_data_27_13;
    assign token_in_vec_13[23] = token_27_13;
    assign in_chan_dep_vld_vec_13[24] = dep_chan_vld_28_13;
    assign in_chan_dep_data_vec_13[999 : 960] = dep_chan_data_28_13;
    assign token_in_vec_13[24] = token_28_13;
    assign in_chan_dep_vld_vec_13[25] = dep_chan_vld_29_13;
    assign in_chan_dep_data_vec_13[1039 : 1000] = dep_chan_data_29_13;
    assign token_in_vec_13[25] = token_29_13;
    assign in_chan_dep_vld_vec_13[26] = dep_chan_vld_30_13;
    assign in_chan_dep_data_vec_13[1079 : 1040] = dep_chan_data_30_13;
    assign token_in_vec_13[26] = token_30_13;
    assign in_chan_dep_vld_vec_13[27] = dep_chan_vld_31_13;
    assign in_chan_dep_data_vec_13[1119 : 1080] = dep_chan_data_31_13;
    assign token_in_vec_13[27] = token_31_13;
    assign in_chan_dep_vld_vec_13[28] = dep_chan_vld_32_13;
    assign in_chan_dep_data_vec_13[1159 : 1120] = dep_chan_data_32_13;
    assign token_in_vec_13[28] = token_32_13;
    assign in_chan_dep_vld_vec_13[29] = dep_chan_vld_33_13;
    assign in_chan_dep_data_vec_13[1199 : 1160] = dep_chan_data_33_13;
    assign token_in_vec_13[29] = token_33_13;
    assign in_chan_dep_vld_vec_13[30] = dep_chan_vld_34_13;
    assign in_chan_dep_data_vec_13[1239 : 1200] = dep_chan_data_34_13;
    assign token_in_vec_13[30] = token_34_13;
    assign in_chan_dep_vld_vec_13[31] = dep_chan_vld_35_13;
    assign in_chan_dep_data_vec_13[1279 : 1240] = dep_chan_data_35_13;
    assign token_in_vec_13[31] = token_35_13;
    assign in_chan_dep_vld_vec_13[32] = dep_chan_vld_36_13;
    assign in_chan_dep_data_vec_13[1319 : 1280] = dep_chan_data_36_13;
    assign token_in_vec_13[32] = token_36_13;
    assign dep_chan_vld_13_12 = out_chan_dep_vld_vec_13[0];
    assign dep_chan_data_13_12 = out_chan_dep_data_13;
    assign token_13_12 = token_out_vec_13[0];
    assign dep_chan_vld_13_14 = out_chan_dep_vld_vec_13[1];
    assign dep_chan_data_13_14 = out_chan_dep_data_13;
    assign token_13_14 = token_out_vec_13[1];
    assign dep_chan_vld_13_0 = out_chan_dep_vld_vec_13[2];
    assign dep_chan_data_13_0 = out_chan_dep_data_13;
    assign token_13_0 = token_out_vec_13[2];
    assign dep_chan_vld_13_1 = out_chan_dep_vld_vec_13[3];
    assign dep_chan_data_13_1 = out_chan_dep_data_13;
    assign token_13_1 = token_out_vec_13[3];
    assign dep_chan_vld_13_3 = out_chan_dep_vld_vec_13[4];
    assign dep_chan_data_13_3 = out_chan_dep_data_13;
    assign token_13_3 = token_out_vec_13[4];
    assign dep_chan_vld_13_6 = out_chan_dep_vld_vec_13[5];
    assign dep_chan_data_13_6 = out_chan_dep_data_13;
    assign token_13_6 = token_out_vec_13[5];
    assign dep_chan_vld_13_7 = out_chan_dep_vld_vec_13[6];
    assign dep_chan_data_13_7 = out_chan_dep_data_13;
    assign token_13_7 = token_out_vec_13[6];
    assign dep_chan_vld_13_8 = out_chan_dep_vld_vec_13[7];
    assign dep_chan_data_13_8 = out_chan_dep_data_13;
    assign token_13_8 = token_out_vec_13[7];
    assign dep_chan_vld_13_9 = out_chan_dep_vld_vec_13[8];
    assign dep_chan_data_13_9 = out_chan_dep_data_13;
    assign token_13_9 = token_out_vec_13[8];
    assign dep_chan_vld_13_10 = out_chan_dep_vld_vec_13[9];
    assign dep_chan_data_13_10 = out_chan_dep_data_13;
    assign token_13_10 = token_out_vec_13[9];
    assign dep_chan_vld_13_11 = out_chan_dep_vld_vec_13[10];
    assign dep_chan_data_13_11 = out_chan_dep_data_13;
    assign token_13_11 = token_out_vec_13[10];
    assign dep_chan_vld_13_15 = out_chan_dep_vld_vec_13[11];
    assign dep_chan_data_13_15 = out_chan_dep_data_13;
    assign token_13_15 = token_out_vec_13[11];
    assign dep_chan_vld_13_16 = out_chan_dep_vld_vec_13[12];
    assign dep_chan_data_13_16 = out_chan_dep_data_13;
    assign token_13_16 = token_out_vec_13[12];
    assign dep_chan_vld_13_17 = out_chan_dep_vld_vec_13[13];
    assign dep_chan_data_13_17 = out_chan_dep_data_13;
    assign token_13_17 = token_out_vec_13[13];
    assign dep_chan_vld_13_18 = out_chan_dep_vld_vec_13[14];
    assign dep_chan_data_13_18 = out_chan_dep_data_13;
    assign token_13_18 = token_out_vec_13[14];
    assign dep_chan_vld_13_19 = out_chan_dep_vld_vec_13[15];
    assign dep_chan_data_13_19 = out_chan_dep_data_13;
    assign token_13_19 = token_out_vec_13[15];
    assign dep_chan_vld_13_20 = out_chan_dep_vld_vec_13[16];
    assign dep_chan_data_13_20 = out_chan_dep_data_13;
    assign token_13_20 = token_out_vec_13[16];
    assign dep_chan_vld_13_21 = out_chan_dep_vld_vec_13[17];
    assign dep_chan_data_13_21 = out_chan_dep_data_13;
    assign token_13_21 = token_out_vec_13[17];
    assign dep_chan_vld_13_22 = out_chan_dep_vld_vec_13[18];
    assign dep_chan_data_13_22 = out_chan_dep_data_13;
    assign token_13_22 = token_out_vec_13[18];
    assign dep_chan_vld_13_23 = out_chan_dep_vld_vec_13[19];
    assign dep_chan_data_13_23 = out_chan_dep_data_13;
    assign token_13_23 = token_out_vec_13[19];
    assign dep_chan_vld_13_24 = out_chan_dep_vld_vec_13[20];
    assign dep_chan_data_13_24 = out_chan_dep_data_13;
    assign token_13_24 = token_out_vec_13[20];
    assign dep_chan_vld_13_25 = out_chan_dep_vld_vec_13[21];
    assign dep_chan_data_13_25 = out_chan_dep_data_13;
    assign token_13_25 = token_out_vec_13[21];
    assign dep_chan_vld_13_26 = out_chan_dep_vld_vec_13[22];
    assign dep_chan_data_13_26 = out_chan_dep_data_13;
    assign token_13_26 = token_out_vec_13[22];
    assign dep_chan_vld_13_27 = out_chan_dep_vld_vec_13[23];
    assign dep_chan_data_13_27 = out_chan_dep_data_13;
    assign token_13_27 = token_out_vec_13[23];
    assign dep_chan_vld_13_28 = out_chan_dep_vld_vec_13[24];
    assign dep_chan_data_13_28 = out_chan_dep_data_13;
    assign token_13_28 = token_out_vec_13[24];
    assign dep_chan_vld_13_29 = out_chan_dep_vld_vec_13[25];
    assign dep_chan_data_13_29 = out_chan_dep_data_13;
    assign token_13_29 = token_out_vec_13[25];
    assign dep_chan_vld_13_30 = out_chan_dep_vld_vec_13[26];
    assign dep_chan_data_13_30 = out_chan_dep_data_13;
    assign token_13_30 = token_out_vec_13[26];
    assign dep_chan_vld_13_31 = out_chan_dep_vld_vec_13[27];
    assign dep_chan_data_13_31 = out_chan_dep_data_13;
    assign token_13_31 = token_out_vec_13[27];
    assign dep_chan_vld_13_32 = out_chan_dep_vld_vec_13[28];
    assign dep_chan_data_13_32 = out_chan_dep_data_13;
    assign token_13_32 = token_out_vec_13[28];
    assign dep_chan_vld_13_33 = out_chan_dep_vld_vec_13[29];
    assign dep_chan_data_13_33 = out_chan_dep_data_13;
    assign token_13_33 = token_out_vec_13[29];
    assign dep_chan_vld_13_34 = out_chan_dep_vld_vec_13[30];
    assign dep_chan_data_13_34 = out_chan_dep_data_13;
    assign token_13_34 = token_out_vec_13[30];
    assign dep_chan_vld_13_35 = out_chan_dep_vld_vec_13[31];
    assign dep_chan_data_13_35 = out_chan_dep_data_13;
    assign token_13_35 = token_out_vec_13[31];
    assign dep_chan_vld_13_36 = out_chan_dep_vld_vec_13[32];
    assign dep_chan_data_13_36 = out_chan_dep_data_13;
    assign token_13_36 = token_out_vec_13[32];

    // Process: ProcessingElement_9_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 14, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_14 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_14),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_14),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_14),
        .token_in_vec(token_in_vec_14),
        .dl_detect_in(dl_detect_out),
        .origin(origin[14]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_14),
        .out_chan_dep_data(out_chan_dep_data_14),
        .token_out_vec(token_out_vec_14),
        .dl_detect_out(dl_in_vec[14]));

    assign proc_14_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_8_blk_n) | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_8_blk_n) | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_WriteC_Flattened_fu_179.cPipes_8_blk_n);
    assign proc_14_data_PIPO_blk[0] = 1'b0;
    assign proc_14_start_FIFO_blk[0] = 1'b0;
    assign proc_14_TLF_FIFO_blk[0] = 1'b0;
    assign proc_14_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_14_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_14[0] = dl_detect_out ? proc_dep_vld_vec_14_reg[0] : (proc_14_data_FIFO_blk[0] | proc_14_data_PIPO_blk[0] | proc_14_start_FIFO_blk[0] | proc_14_TLF_FIFO_blk[0] | proc_14_input_sync_blk[0] | proc_14_output_sync_blk[0]);
    assign proc_14_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_9_blk_n) | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_9_blk_n) | (~ProcessingElement_9_U0.grp_ProcessingElement_9_Pipeline_WriteC_Flattened_fu_179.cPipes_9_blk_n);
    assign proc_14_data_PIPO_blk[1] = 1'b0;
    assign proc_14_start_FIFO_blk[1] = 1'b0;
    assign proc_14_TLF_FIFO_blk[1] = 1'b0;
    assign proc_14_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_14_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_14[1] = dl_detect_out ? proc_dep_vld_vec_14_reg[1] : (proc_14_data_FIFO_blk[1] | proc_14_data_PIPO_blk[1] | proc_14_start_FIFO_blk[1] | proc_14_TLF_FIFO_blk[1] | proc_14_input_sync_blk[1] | proc_14_output_sync_blk[1]);
    assign proc_14_data_FIFO_blk[2] = 1'b0;
    assign proc_14_data_PIPO_blk[2] = 1'b0;
    assign proc_14_start_FIFO_blk[2] = 1'b0;
    assign proc_14_TLF_FIFO_blk[2] = 1'b0;
    assign proc_14_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_14_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_14[2] = dl_detect_out ? proc_dep_vld_vec_14_reg[2] : (proc_14_data_FIFO_blk[2] | proc_14_data_PIPO_blk[2] | proc_14_start_FIFO_blk[2] | proc_14_TLF_FIFO_blk[2] | proc_14_input_sync_blk[2] | proc_14_output_sync_blk[2]);
    assign proc_14_data_FIFO_blk[3] = 1'b0;
    assign proc_14_data_PIPO_blk[3] = 1'b0;
    assign proc_14_start_FIFO_blk[3] = 1'b0;
    assign proc_14_TLF_FIFO_blk[3] = 1'b0;
    assign proc_14_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_14_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_14[3] = dl_detect_out ? proc_dep_vld_vec_14_reg[3] : (proc_14_data_FIFO_blk[3] | proc_14_data_PIPO_blk[3] | proc_14_start_FIFO_blk[3] | proc_14_TLF_FIFO_blk[3] | proc_14_input_sync_blk[3] | proc_14_output_sync_blk[3]);
    assign proc_14_data_FIFO_blk[4] = 1'b0;
    assign proc_14_data_PIPO_blk[4] = 1'b0;
    assign proc_14_start_FIFO_blk[4] = 1'b0;
    assign proc_14_TLF_FIFO_blk[4] = 1'b0;
    assign proc_14_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_14_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_14[4] = dl_detect_out ? proc_dep_vld_vec_14_reg[4] : (proc_14_data_FIFO_blk[4] | proc_14_data_PIPO_blk[4] | proc_14_start_FIFO_blk[4] | proc_14_TLF_FIFO_blk[4] | proc_14_input_sync_blk[4] | proc_14_output_sync_blk[4]);
    assign proc_14_data_FIFO_blk[5] = 1'b0;
    assign proc_14_data_PIPO_blk[5] = 1'b0;
    assign proc_14_start_FIFO_blk[5] = 1'b0;
    assign proc_14_TLF_FIFO_blk[5] = 1'b0;
    assign proc_14_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_14_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_14[5] = dl_detect_out ? proc_dep_vld_vec_14_reg[5] : (proc_14_data_FIFO_blk[5] | proc_14_data_PIPO_blk[5] | proc_14_start_FIFO_blk[5] | proc_14_TLF_FIFO_blk[5] | proc_14_input_sync_blk[5] | proc_14_output_sync_blk[5]);
    assign proc_14_data_FIFO_blk[6] = 1'b0;
    assign proc_14_data_PIPO_blk[6] = 1'b0;
    assign proc_14_start_FIFO_blk[6] = 1'b0;
    assign proc_14_TLF_FIFO_blk[6] = 1'b0;
    assign proc_14_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_14_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_14[6] = dl_detect_out ? proc_dep_vld_vec_14_reg[6] : (proc_14_data_FIFO_blk[6] | proc_14_data_PIPO_blk[6] | proc_14_start_FIFO_blk[6] | proc_14_TLF_FIFO_blk[6] | proc_14_input_sync_blk[6] | proc_14_output_sync_blk[6]);
    assign proc_14_data_FIFO_blk[7] = 1'b0;
    assign proc_14_data_PIPO_blk[7] = 1'b0;
    assign proc_14_start_FIFO_blk[7] = 1'b0;
    assign proc_14_TLF_FIFO_blk[7] = 1'b0;
    assign proc_14_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_14_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_14[7] = dl_detect_out ? proc_dep_vld_vec_14_reg[7] : (proc_14_data_FIFO_blk[7] | proc_14_data_PIPO_blk[7] | proc_14_start_FIFO_blk[7] | proc_14_TLF_FIFO_blk[7] | proc_14_input_sync_blk[7] | proc_14_output_sync_blk[7]);
    assign proc_14_data_FIFO_blk[8] = 1'b0;
    assign proc_14_data_PIPO_blk[8] = 1'b0;
    assign proc_14_start_FIFO_blk[8] = 1'b0;
    assign proc_14_TLF_FIFO_blk[8] = 1'b0;
    assign proc_14_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_14_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_14[8] = dl_detect_out ? proc_dep_vld_vec_14_reg[8] : (proc_14_data_FIFO_blk[8] | proc_14_data_PIPO_blk[8] | proc_14_start_FIFO_blk[8] | proc_14_TLF_FIFO_blk[8] | proc_14_input_sync_blk[8] | proc_14_output_sync_blk[8]);
    assign proc_14_data_FIFO_blk[9] = 1'b0;
    assign proc_14_data_PIPO_blk[9] = 1'b0;
    assign proc_14_start_FIFO_blk[9] = 1'b0;
    assign proc_14_TLF_FIFO_blk[9] = 1'b0;
    assign proc_14_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_14_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_14[9] = dl_detect_out ? proc_dep_vld_vec_14_reg[9] : (proc_14_data_FIFO_blk[9] | proc_14_data_PIPO_blk[9] | proc_14_start_FIFO_blk[9] | proc_14_TLF_FIFO_blk[9] | proc_14_input_sync_blk[9] | proc_14_output_sync_blk[9]);
    assign proc_14_data_FIFO_blk[10] = 1'b0;
    assign proc_14_data_PIPO_blk[10] = 1'b0;
    assign proc_14_start_FIFO_blk[10] = 1'b0;
    assign proc_14_TLF_FIFO_blk[10] = 1'b0;
    assign proc_14_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_14_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_14[10] = dl_detect_out ? proc_dep_vld_vec_14_reg[10] : (proc_14_data_FIFO_blk[10] | proc_14_data_PIPO_blk[10] | proc_14_start_FIFO_blk[10] | proc_14_TLF_FIFO_blk[10] | proc_14_input_sync_blk[10] | proc_14_output_sync_blk[10]);
    assign proc_14_data_FIFO_blk[11] = 1'b0;
    assign proc_14_data_PIPO_blk[11] = 1'b0;
    assign proc_14_start_FIFO_blk[11] = 1'b0;
    assign proc_14_TLF_FIFO_blk[11] = 1'b0;
    assign proc_14_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_14_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_14[11] = dl_detect_out ? proc_dep_vld_vec_14_reg[11] : (proc_14_data_FIFO_blk[11] | proc_14_data_PIPO_blk[11] | proc_14_start_FIFO_blk[11] | proc_14_TLF_FIFO_blk[11] | proc_14_input_sync_blk[11] | proc_14_output_sync_blk[11]);
    assign proc_14_data_FIFO_blk[12] = 1'b0;
    assign proc_14_data_PIPO_blk[12] = 1'b0;
    assign proc_14_start_FIFO_blk[12] = 1'b0;
    assign proc_14_TLF_FIFO_blk[12] = 1'b0;
    assign proc_14_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_14_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_14[12] = dl_detect_out ? proc_dep_vld_vec_14_reg[12] : (proc_14_data_FIFO_blk[12] | proc_14_data_PIPO_blk[12] | proc_14_start_FIFO_blk[12] | proc_14_TLF_FIFO_blk[12] | proc_14_input_sync_blk[12] | proc_14_output_sync_blk[12]);
    assign proc_14_data_FIFO_blk[13] = 1'b0;
    assign proc_14_data_PIPO_blk[13] = 1'b0;
    assign proc_14_start_FIFO_blk[13] = 1'b0;
    assign proc_14_TLF_FIFO_blk[13] = 1'b0;
    assign proc_14_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_14_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_14[13] = dl_detect_out ? proc_dep_vld_vec_14_reg[13] : (proc_14_data_FIFO_blk[13] | proc_14_data_PIPO_blk[13] | proc_14_start_FIFO_blk[13] | proc_14_TLF_FIFO_blk[13] | proc_14_input_sync_blk[13] | proc_14_output_sync_blk[13]);
    assign proc_14_data_FIFO_blk[14] = 1'b0;
    assign proc_14_data_PIPO_blk[14] = 1'b0;
    assign proc_14_start_FIFO_blk[14] = 1'b0;
    assign proc_14_TLF_FIFO_blk[14] = 1'b0;
    assign proc_14_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_14_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_14[14] = dl_detect_out ? proc_dep_vld_vec_14_reg[14] : (proc_14_data_FIFO_blk[14] | proc_14_data_PIPO_blk[14] | proc_14_start_FIFO_blk[14] | proc_14_TLF_FIFO_blk[14] | proc_14_input_sync_blk[14] | proc_14_output_sync_blk[14]);
    assign proc_14_data_FIFO_blk[15] = 1'b0;
    assign proc_14_data_PIPO_blk[15] = 1'b0;
    assign proc_14_start_FIFO_blk[15] = 1'b0;
    assign proc_14_TLF_FIFO_blk[15] = 1'b0;
    assign proc_14_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_14_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_14[15] = dl_detect_out ? proc_dep_vld_vec_14_reg[15] : (proc_14_data_FIFO_blk[15] | proc_14_data_PIPO_blk[15] | proc_14_start_FIFO_blk[15] | proc_14_TLF_FIFO_blk[15] | proc_14_input_sync_blk[15] | proc_14_output_sync_blk[15]);
    assign proc_14_data_FIFO_blk[16] = 1'b0;
    assign proc_14_data_PIPO_blk[16] = 1'b0;
    assign proc_14_start_FIFO_blk[16] = 1'b0;
    assign proc_14_TLF_FIFO_blk[16] = 1'b0;
    assign proc_14_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_14_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_14[16] = dl_detect_out ? proc_dep_vld_vec_14_reg[16] : (proc_14_data_FIFO_blk[16] | proc_14_data_PIPO_blk[16] | proc_14_start_FIFO_blk[16] | proc_14_TLF_FIFO_blk[16] | proc_14_input_sync_blk[16] | proc_14_output_sync_blk[16]);
    assign proc_14_data_FIFO_blk[17] = 1'b0;
    assign proc_14_data_PIPO_blk[17] = 1'b0;
    assign proc_14_start_FIFO_blk[17] = 1'b0;
    assign proc_14_TLF_FIFO_blk[17] = 1'b0;
    assign proc_14_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_14_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_14[17] = dl_detect_out ? proc_dep_vld_vec_14_reg[17] : (proc_14_data_FIFO_blk[17] | proc_14_data_PIPO_blk[17] | proc_14_start_FIFO_blk[17] | proc_14_TLF_FIFO_blk[17] | proc_14_input_sync_blk[17] | proc_14_output_sync_blk[17]);
    assign proc_14_data_FIFO_blk[18] = 1'b0;
    assign proc_14_data_PIPO_blk[18] = 1'b0;
    assign proc_14_start_FIFO_blk[18] = 1'b0;
    assign proc_14_TLF_FIFO_blk[18] = 1'b0;
    assign proc_14_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_14_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_14[18] = dl_detect_out ? proc_dep_vld_vec_14_reg[18] : (proc_14_data_FIFO_blk[18] | proc_14_data_PIPO_blk[18] | proc_14_start_FIFO_blk[18] | proc_14_TLF_FIFO_blk[18] | proc_14_input_sync_blk[18] | proc_14_output_sync_blk[18]);
    assign proc_14_data_FIFO_blk[19] = 1'b0;
    assign proc_14_data_PIPO_blk[19] = 1'b0;
    assign proc_14_start_FIFO_blk[19] = 1'b0;
    assign proc_14_TLF_FIFO_blk[19] = 1'b0;
    assign proc_14_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_14_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_14[19] = dl_detect_out ? proc_dep_vld_vec_14_reg[19] : (proc_14_data_FIFO_blk[19] | proc_14_data_PIPO_blk[19] | proc_14_start_FIFO_blk[19] | proc_14_TLF_FIFO_blk[19] | proc_14_input_sync_blk[19] | proc_14_output_sync_blk[19]);
    assign proc_14_data_FIFO_blk[20] = 1'b0;
    assign proc_14_data_PIPO_blk[20] = 1'b0;
    assign proc_14_start_FIFO_blk[20] = 1'b0;
    assign proc_14_TLF_FIFO_blk[20] = 1'b0;
    assign proc_14_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_14_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_14[20] = dl_detect_out ? proc_dep_vld_vec_14_reg[20] : (proc_14_data_FIFO_blk[20] | proc_14_data_PIPO_blk[20] | proc_14_start_FIFO_blk[20] | proc_14_TLF_FIFO_blk[20] | proc_14_input_sync_blk[20] | proc_14_output_sync_blk[20]);
    assign proc_14_data_FIFO_blk[21] = 1'b0;
    assign proc_14_data_PIPO_blk[21] = 1'b0;
    assign proc_14_start_FIFO_blk[21] = 1'b0;
    assign proc_14_TLF_FIFO_blk[21] = 1'b0;
    assign proc_14_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_14_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_14[21] = dl_detect_out ? proc_dep_vld_vec_14_reg[21] : (proc_14_data_FIFO_blk[21] | proc_14_data_PIPO_blk[21] | proc_14_start_FIFO_blk[21] | proc_14_TLF_FIFO_blk[21] | proc_14_input_sync_blk[21] | proc_14_output_sync_blk[21]);
    assign proc_14_data_FIFO_blk[22] = 1'b0;
    assign proc_14_data_PIPO_blk[22] = 1'b0;
    assign proc_14_start_FIFO_blk[22] = 1'b0;
    assign proc_14_TLF_FIFO_blk[22] = 1'b0;
    assign proc_14_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_14_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_14[22] = dl_detect_out ? proc_dep_vld_vec_14_reg[22] : (proc_14_data_FIFO_blk[22] | proc_14_data_PIPO_blk[22] | proc_14_start_FIFO_blk[22] | proc_14_TLF_FIFO_blk[22] | proc_14_input_sync_blk[22] | proc_14_output_sync_blk[22]);
    assign proc_14_data_FIFO_blk[23] = 1'b0;
    assign proc_14_data_PIPO_blk[23] = 1'b0;
    assign proc_14_start_FIFO_blk[23] = 1'b0;
    assign proc_14_TLF_FIFO_blk[23] = 1'b0;
    assign proc_14_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_14_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_14[23] = dl_detect_out ? proc_dep_vld_vec_14_reg[23] : (proc_14_data_FIFO_blk[23] | proc_14_data_PIPO_blk[23] | proc_14_start_FIFO_blk[23] | proc_14_TLF_FIFO_blk[23] | proc_14_input_sync_blk[23] | proc_14_output_sync_blk[23]);
    assign proc_14_data_FIFO_blk[24] = 1'b0;
    assign proc_14_data_PIPO_blk[24] = 1'b0;
    assign proc_14_start_FIFO_blk[24] = 1'b0;
    assign proc_14_TLF_FIFO_blk[24] = 1'b0;
    assign proc_14_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_14_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_14[24] = dl_detect_out ? proc_dep_vld_vec_14_reg[24] : (proc_14_data_FIFO_blk[24] | proc_14_data_PIPO_blk[24] | proc_14_start_FIFO_blk[24] | proc_14_TLF_FIFO_blk[24] | proc_14_input_sync_blk[24] | proc_14_output_sync_blk[24]);
    assign proc_14_data_FIFO_blk[25] = 1'b0;
    assign proc_14_data_PIPO_blk[25] = 1'b0;
    assign proc_14_start_FIFO_blk[25] = 1'b0;
    assign proc_14_TLF_FIFO_blk[25] = 1'b0;
    assign proc_14_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_14_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_14[25] = dl_detect_out ? proc_dep_vld_vec_14_reg[25] : (proc_14_data_FIFO_blk[25] | proc_14_data_PIPO_blk[25] | proc_14_start_FIFO_blk[25] | proc_14_TLF_FIFO_blk[25] | proc_14_input_sync_blk[25] | proc_14_output_sync_blk[25]);
    assign proc_14_data_FIFO_blk[26] = 1'b0;
    assign proc_14_data_PIPO_blk[26] = 1'b0;
    assign proc_14_start_FIFO_blk[26] = 1'b0;
    assign proc_14_TLF_FIFO_blk[26] = 1'b0;
    assign proc_14_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_14_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_14[26] = dl_detect_out ? proc_dep_vld_vec_14_reg[26] : (proc_14_data_FIFO_blk[26] | proc_14_data_PIPO_blk[26] | proc_14_start_FIFO_blk[26] | proc_14_TLF_FIFO_blk[26] | proc_14_input_sync_blk[26] | proc_14_output_sync_blk[26]);
    assign proc_14_data_FIFO_blk[27] = 1'b0;
    assign proc_14_data_PIPO_blk[27] = 1'b0;
    assign proc_14_start_FIFO_blk[27] = 1'b0;
    assign proc_14_TLF_FIFO_blk[27] = 1'b0;
    assign proc_14_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_14_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_14[27] = dl_detect_out ? proc_dep_vld_vec_14_reg[27] : (proc_14_data_FIFO_blk[27] | proc_14_data_PIPO_blk[27] | proc_14_start_FIFO_blk[27] | proc_14_TLF_FIFO_blk[27] | proc_14_input_sync_blk[27] | proc_14_output_sync_blk[27]);
    assign proc_14_data_FIFO_blk[28] = 1'b0;
    assign proc_14_data_PIPO_blk[28] = 1'b0;
    assign proc_14_start_FIFO_blk[28] = 1'b0;
    assign proc_14_TLF_FIFO_blk[28] = 1'b0;
    assign proc_14_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_14_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_14[28] = dl_detect_out ? proc_dep_vld_vec_14_reg[28] : (proc_14_data_FIFO_blk[28] | proc_14_data_PIPO_blk[28] | proc_14_start_FIFO_blk[28] | proc_14_TLF_FIFO_blk[28] | proc_14_input_sync_blk[28] | proc_14_output_sync_blk[28]);
    assign proc_14_data_FIFO_blk[29] = 1'b0;
    assign proc_14_data_PIPO_blk[29] = 1'b0;
    assign proc_14_start_FIFO_blk[29] = 1'b0;
    assign proc_14_TLF_FIFO_blk[29] = 1'b0;
    assign proc_14_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_14_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_14[29] = dl_detect_out ? proc_dep_vld_vec_14_reg[29] : (proc_14_data_FIFO_blk[29] | proc_14_data_PIPO_blk[29] | proc_14_start_FIFO_blk[29] | proc_14_TLF_FIFO_blk[29] | proc_14_input_sync_blk[29] | proc_14_output_sync_blk[29]);
    assign proc_14_data_FIFO_blk[30] = 1'b0;
    assign proc_14_data_PIPO_blk[30] = 1'b0;
    assign proc_14_start_FIFO_blk[30] = 1'b0;
    assign proc_14_TLF_FIFO_blk[30] = 1'b0;
    assign proc_14_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_14_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_14[30] = dl_detect_out ? proc_dep_vld_vec_14_reg[30] : (proc_14_data_FIFO_blk[30] | proc_14_data_PIPO_blk[30] | proc_14_start_FIFO_blk[30] | proc_14_TLF_FIFO_blk[30] | proc_14_input_sync_blk[30] | proc_14_output_sync_blk[30]);
    assign proc_14_data_FIFO_blk[31] = 1'b0;
    assign proc_14_data_PIPO_blk[31] = 1'b0;
    assign proc_14_start_FIFO_blk[31] = 1'b0;
    assign proc_14_TLF_FIFO_blk[31] = 1'b0;
    assign proc_14_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_14_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_14[31] = dl_detect_out ? proc_dep_vld_vec_14_reg[31] : (proc_14_data_FIFO_blk[31] | proc_14_data_PIPO_blk[31] | proc_14_start_FIFO_blk[31] | proc_14_TLF_FIFO_blk[31] | proc_14_input_sync_blk[31] | proc_14_output_sync_blk[31]);
    assign proc_14_data_FIFO_blk[32] = 1'b0;
    assign proc_14_data_PIPO_blk[32] = 1'b0;
    assign proc_14_start_FIFO_blk[32] = 1'b0;
    assign proc_14_TLF_FIFO_blk[32] = 1'b0;
    assign proc_14_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_9_U0_ap_ready & ProcessingElement_9_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_14_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_14[32] = dl_detect_out ? proc_dep_vld_vec_14_reg[32] : (proc_14_data_FIFO_blk[32] | proc_14_data_PIPO_blk[32] | proc_14_start_FIFO_blk[32] | proc_14_TLF_FIFO_blk[32] | proc_14_input_sync_blk[32] | proc_14_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_14_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_14_reg <= proc_dep_vld_vec_14;
        end
    end
    assign in_chan_dep_vld_vec_14[0] = dep_chan_vld_0_14;
    assign in_chan_dep_data_vec_14[39 : 0] = dep_chan_data_0_14;
    assign token_in_vec_14[0] = token_0_14;
    assign in_chan_dep_vld_vec_14[1] = dep_chan_vld_1_14;
    assign in_chan_dep_data_vec_14[79 : 40] = dep_chan_data_1_14;
    assign token_in_vec_14[1] = token_1_14;
    assign in_chan_dep_vld_vec_14[2] = dep_chan_vld_3_14;
    assign in_chan_dep_data_vec_14[119 : 80] = dep_chan_data_3_14;
    assign token_in_vec_14[2] = token_3_14;
    assign in_chan_dep_vld_vec_14[3] = dep_chan_vld_6_14;
    assign in_chan_dep_data_vec_14[159 : 120] = dep_chan_data_6_14;
    assign token_in_vec_14[3] = token_6_14;
    assign in_chan_dep_vld_vec_14[4] = dep_chan_vld_7_14;
    assign in_chan_dep_data_vec_14[199 : 160] = dep_chan_data_7_14;
    assign token_in_vec_14[4] = token_7_14;
    assign in_chan_dep_vld_vec_14[5] = dep_chan_vld_8_14;
    assign in_chan_dep_data_vec_14[239 : 200] = dep_chan_data_8_14;
    assign token_in_vec_14[5] = token_8_14;
    assign in_chan_dep_vld_vec_14[6] = dep_chan_vld_9_14;
    assign in_chan_dep_data_vec_14[279 : 240] = dep_chan_data_9_14;
    assign token_in_vec_14[6] = token_9_14;
    assign in_chan_dep_vld_vec_14[7] = dep_chan_vld_10_14;
    assign in_chan_dep_data_vec_14[319 : 280] = dep_chan_data_10_14;
    assign token_in_vec_14[7] = token_10_14;
    assign in_chan_dep_vld_vec_14[8] = dep_chan_vld_11_14;
    assign in_chan_dep_data_vec_14[359 : 320] = dep_chan_data_11_14;
    assign token_in_vec_14[8] = token_11_14;
    assign in_chan_dep_vld_vec_14[9] = dep_chan_vld_12_14;
    assign in_chan_dep_data_vec_14[399 : 360] = dep_chan_data_12_14;
    assign token_in_vec_14[9] = token_12_14;
    assign in_chan_dep_vld_vec_14[10] = dep_chan_vld_13_14;
    assign in_chan_dep_data_vec_14[439 : 400] = dep_chan_data_13_14;
    assign token_in_vec_14[10] = token_13_14;
    assign in_chan_dep_vld_vec_14[11] = dep_chan_vld_15_14;
    assign in_chan_dep_data_vec_14[479 : 440] = dep_chan_data_15_14;
    assign token_in_vec_14[11] = token_15_14;
    assign in_chan_dep_vld_vec_14[12] = dep_chan_vld_16_14;
    assign in_chan_dep_data_vec_14[519 : 480] = dep_chan_data_16_14;
    assign token_in_vec_14[12] = token_16_14;
    assign in_chan_dep_vld_vec_14[13] = dep_chan_vld_17_14;
    assign in_chan_dep_data_vec_14[559 : 520] = dep_chan_data_17_14;
    assign token_in_vec_14[13] = token_17_14;
    assign in_chan_dep_vld_vec_14[14] = dep_chan_vld_18_14;
    assign in_chan_dep_data_vec_14[599 : 560] = dep_chan_data_18_14;
    assign token_in_vec_14[14] = token_18_14;
    assign in_chan_dep_vld_vec_14[15] = dep_chan_vld_19_14;
    assign in_chan_dep_data_vec_14[639 : 600] = dep_chan_data_19_14;
    assign token_in_vec_14[15] = token_19_14;
    assign in_chan_dep_vld_vec_14[16] = dep_chan_vld_20_14;
    assign in_chan_dep_data_vec_14[679 : 640] = dep_chan_data_20_14;
    assign token_in_vec_14[16] = token_20_14;
    assign in_chan_dep_vld_vec_14[17] = dep_chan_vld_21_14;
    assign in_chan_dep_data_vec_14[719 : 680] = dep_chan_data_21_14;
    assign token_in_vec_14[17] = token_21_14;
    assign in_chan_dep_vld_vec_14[18] = dep_chan_vld_22_14;
    assign in_chan_dep_data_vec_14[759 : 720] = dep_chan_data_22_14;
    assign token_in_vec_14[18] = token_22_14;
    assign in_chan_dep_vld_vec_14[19] = dep_chan_vld_23_14;
    assign in_chan_dep_data_vec_14[799 : 760] = dep_chan_data_23_14;
    assign token_in_vec_14[19] = token_23_14;
    assign in_chan_dep_vld_vec_14[20] = dep_chan_vld_24_14;
    assign in_chan_dep_data_vec_14[839 : 800] = dep_chan_data_24_14;
    assign token_in_vec_14[20] = token_24_14;
    assign in_chan_dep_vld_vec_14[21] = dep_chan_vld_25_14;
    assign in_chan_dep_data_vec_14[879 : 840] = dep_chan_data_25_14;
    assign token_in_vec_14[21] = token_25_14;
    assign in_chan_dep_vld_vec_14[22] = dep_chan_vld_26_14;
    assign in_chan_dep_data_vec_14[919 : 880] = dep_chan_data_26_14;
    assign token_in_vec_14[22] = token_26_14;
    assign in_chan_dep_vld_vec_14[23] = dep_chan_vld_27_14;
    assign in_chan_dep_data_vec_14[959 : 920] = dep_chan_data_27_14;
    assign token_in_vec_14[23] = token_27_14;
    assign in_chan_dep_vld_vec_14[24] = dep_chan_vld_28_14;
    assign in_chan_dep_data_vec_14[999 : 960] = dep_chan_data_28_14;
    assign token_in_vec_14[24] = token_28_14;
    assign in_chan_dep_vld_vec_14[25] = dep_chan_vld_29_14;
    assign in_chan_dep_data_vec_14[1039 : 1000] = dep_chan_data_29_14;
    assign token_in_vec_14[25] = token_29_14;
    assign in_chan_dep_vld_vec_14[26] = dep_chan_vld_30_14;
    assign in_chan_dep_data_vec_14[1079 : 1040] = dep_chan_data_30_14;
    assign token_in_vec_14[26] = token_30_14;
    assign in_chan_dep_vld_vec_14[27] = dep_chan_vld_31_14;
    assign in_chan_dep_data_vec_14[1119 : 1080] = dep_chan_data_31_14;
    assign token_in_vec_14[27] = token_31_14;
    assign in_chan_dep_vld_vec_14[28] = dep_chan_vld_32_14;
    assign in_chan_dep_data_vec_14[1159 : 1120] = dep_chan_data_32_14;
    assign token_in_vec_14[28] = token_32_14;
    assign in_chan_dep_vld_vec_14[29] = dep_chan_vld_33_14;
    assign in_chan_dep_data_vec_14[1199 : 1160] = dep_chan_data_33_14;
    assign token_in_vec_14[29] = token_33_14;
    assign in_chan_dep_vld_vec_14[30] = dep_chan_vld_34_14;
    assign in_chan_dep_data_vec_14[1239 : 1200] = dep_chan_data_34_14;
    assign token_in_vec_14[30] = token_34_14;
    assign in_chan_dep_vld_vec_14[31] = dep_chan_vld_35_14;
    assign in_chan_dep_data_vec_14[1279 : 1240] = dep_chan_data_35_14;
    assign token_in_vec_14[31] = token_35_14;
    assign in_chan_dep_vld_vec_14[32] = dep_chan_vld_36_14;
    assign in_chan_dep_data_vec_14[1319 : 1280] = dep_chan_data_36_14;
    assign token_in_vec_14[32] = token_36_14;
    assign dep_chan_vld_14_13 = out_chan_dep_vld_vec_14[0];
    assign dep_chan_data_14_13 = out_chan_dep_data_14;
    assign token_14_13 = token_out_vec_14[0];
    assign dep_chan_vld_14_15 = out_chan_dep_vld_vec_14[1];
    assign dep_chan_data_14_15 = out_chan_dep_data_14;
    assign token_14_15 = token_out_vec_14[1];
    assign dep_chan_vld_14_0 = out_chan_dep_vld_vec_14[2];
    assign dep_chan_data_14_0 = out_chan_dep_data_14;
    assign token_14_0 = token_out_vec_14[2];
    assign dep_chan_vld_14_1 = out_chan_dep_vld_vec_14[3];
    assign dep_chan_data_14_1 = out_chan_dep_data_14;
    assign token_14_1 = token_out_vec_14[3];
    assign dep_chan_vld_14_3 = out_chan_dep_vld_vec_14[4];
    assign dep_chan_data_14_3 = out_chan_dep_data_14;
    assign token_14_3 = token_out_vec_14[4];
    assign dep_chan_vld_14_6 = out_chan_dep_vld_vec_14[5];
    assign dep_chan_data_14_6 = out_chan_dep_data_14;
    assign token_14_6 = token_out_vec_14[5];
    assign dep_chan_vld_14_7 = out_chan_dep_vld_vec_14[6];
    assign dep_chan_data_14_7 = out_chan_dep_data_14;
    assign token_14_7 = token_out_vec_14[6];
    assign dep_chan_vld_14_8 = out_chan_dep_vld_vec_14[7];
    assign dep_chan_data_14_8 = out_chan_dep_data_14;
    assign token_14_8 = token_out_vec_14[7];
    assign dep_chan_vld_14_9 = out_chan_dep_vld_vec_14[8];
    assign dep_chan_data_14_9 = out_chan_dep_data_14;
    assign token_14_9 = token_out_vec_14[8];
    assign dep_chan_vld_14_10 = out_chan_dep_vld_vec_14[9];
    assign dep_chan_data_14_10 = out_chan_dep_data_14;
    assign token_14_10 = token_out_vec_14[9];
    assign dep_chan_vld_14_11 = out_chan_dep_vld_vec_14[10];
    assign dep_chan_data_14_11 = out_chan_dep_data_14;
    assign token_14_11 = token_out_vec_14[10];
    assign dep_chan_vld_14_12 = out_chan_dep_vld_vec_14[11];
    assign dep_chan_data_14_12 = out_chan_dep_data_14;
    assign token_14_12 = token_out_vec_14[11];
    assign dep_chan_vld_14_16 = out_chan_dep_vld_vec_14[12];
    assign dep_chan_data_14_16 = out_chan_dep_data_14;
    assign token_14_16 = token_out_vec_14[12];
    assign dep_chan_vld_14_17 = out_chan_dep_vld_vec_14[13];
    assign dep_chan_data_14_17 = out_chan_dep_data_14;
    assign token_14_17 = token_out_vec_14[13];
    assign dep_chan_vld_14_18 = out_chan_dep_vld_vec_14[14];
    assign dep_chan_data_14_18 = out_chan_dep_data_14;
    assign token_14_18 = token_out_vec_14[14];
    assign dep_chan_vld_14_19 = out_chan_dep_vld_vec_14[15];
    assign dep_chan_data_14_19 = out_chan_dep_data_14;
    assign token_14_19 = token_out_vec_14[15];
    assign dep_chan_vld_14_20 = out_chan_dep_vld_vec_14[16];
    assign dep_chan_data_14_20 = out_chan_dep_data_14;
    assign token_14_20 = token_out_vec_14[16];
    assign dep_chan_vld_14_21 = out_chan_dep_vld_vec_14[17];
    assign dep_chan_data_14_21 = out_chan_dep_data_14;
    assign token_14_21 = token_out_vec_14[17];
    assign dep_chan_vld_14_22 = out_chan_dep_vld_vec_14[18];
    assign dep_chan_data_14_22 = out_chan_dep_data_14;
    assign token_14_22 = token_out_vec_14[18];
    assign dep_chan_vld_14_23 = out_chan_dep_vld_vec_14[19];
    assign dep_chan_data_14_23 = out_chan_dep_data_14;
    assign token_14_23 = token_out_vec_14[19];
    assign dep_chan_vld_14_24 = out_chan_dep_vld_vec_14[20];
    assign dep_chan_data_14_24 = out_chan_dep_data_14;
    assign token_14_24 = token_out_vec_14[20];
    assign dep_chan_vld_14_25 = out_chan_dep_vld_vec_14[21];
    assign dep_chan_data_14_25 = out_chan_dep_data_14;
    assign token_14_25 = token_out_vec_14[21];
    assign dep_chan_vld_14_26 = out_chan_dep_vld_vec_14[22];
    assign dep_chan_data_14_26 = out_chan_dep_data_14;
    assign token_14_26 = token_out_vec_14[22];
    assign dep_chan_vld_14_27 = out_chan_dep_vld_vec_14[23];
    assign dep_chan_data_14_27 = out_chan_dep_data_14;
    assign token_14_27 = token_out_vec_14[23];
    assign dep_chan_vld_14_28 = out_chan_dep_vld_vec_14[24];
    assign dep_chan_data_14_28 = out_chan_dep_data_14;
    assign token_14_28 = token_out_vec_14[24];
    assign dep_chan_vld_14_29 = out_chan_dep_vld_vec_14[25];
    assign dep_chan_data_14_29 = out_chan_dep_data_14;
    assign token_14_29 = token_out_vec_14[25];
    assign dep_chan_vld_14_30 = out_chan_dep_vld_vec_14[26];
    assign dep_chan_data_14_30 = out_chan_dep_data_14;
    assign token_14_30 = token_out_vec_14[26];
    assign dep_chan_vld_14_31 = out_chan_dep_vld_vec_14[27];
    assign dep_chan_data_14_31 = out_chan_dep_data_14;
    assign token_14_31 = token_out_vec_14[27];
    assign dep_chan_vld_14_32 = out_chan_dep_vld_vec_14[28];
    assign dep_chan_data_14_32 = out_chan_dep_data_14;
    assign token_14_32 = token_out_vec_14[28];
    assign dep_chan_vld_14_33 = out_chan_dep_vld_vec_14[29];
    assign dep_chan_data_14_33 = out_chan_dep_data_14;
    assign token_14_33 = token_out_vec_14[29];
    assign dep_chan_vld_14_34 = out_chan_dep_vld_vec_14[30];
    assign dep_chan_data_14_34 = out_chan_dep_data_14;
    assign token_14_34 = token_out_vec_14[30];
    assign dep_chan_vld_14_35 = out_chan_dep_vld_vec_14[31];
    assign dep_chan_data_14_35 = out_chan_dep_data_14;
    assign token_14_35 = token_out_vec_14[31];
    assign dep_chan_vld_14_36 = out_chan_dep_vld_vec_14[32];
    assign dep_chan_data_14_36 = out_chan_dep_data_14;
    assign token_14_36 = token_out_vec_14[32];

    // Process: ProcessingElement_10_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 15, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_15 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_15),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_15),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_15),
        .token_in_vec(token_in_vec_15),
        .dl_detect_in(dl_detect_out),
        .origin(origin[15]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_15),
        .out_chan_dep_data(out_chan_dep_data_15),
        .token_out_vec(token_out_vec_15),
        .dl_detect_out(dl_in_vec[15]));

    assign proc_15_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_9_blk_n) | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_9_blk_n) | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_WriteC_Flattened_fu_179.cPipes_9_blk_n);
    assign proc_15_data_PIPO_blk[0] = 1'b0;
    assign proc_15_start_FIFO_blk[0] = 1'b0;
    assign proc_15_TLF_FIFO_blk[0] = 1'b0;
    assign proc_15_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_15_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_15[0] = dl_detect_out ? proc_dep_vld_vec_15_reg[0] : (proc_15_data_FIFO_blk[0] | proc_15_data_PIPO_blk[0] | proc_15_start_FIFO_blk[0] | proc_15_TLF_FIFO_blk[0] | proc_15_input_sync_blk[0] | proc_15_output_sync_blk[0]);
    assign proc_15_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_10_blk_n) | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_10_blk_n) | (~ProcessingElement_10_U0.grp_ProcessingElement_10_Pipeline_WriteC_Flattened_fu_179.cPipes_10_blk_n);
    assign proc_15_data_PIPO_blk[1] = 1'b0;
    assign proc_15_start_FIFO_blk[1] = 1'b0;
    assign proc_15_TLF_FIFO_blk[1] = 1'b0;
    assign proc_15_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_15_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_15[1] = dl_detect_out ? proc_dep_vld_vec_15_reg[1] : (proc_15_data_FIFO_blk[1] | proc_15_data_PIPO_blk[1] | proc_15_start_FIFO_blk[1] | proc_15_TLF_FIFO_blk[1] | proc_15_input_sync_blk[1] | proc_15_output_sync_blk[1]);
    assign proc_15_data_FIFO_blk[2] = 1'b0;
    assign proc_15_data_PIPO_blk[2] = 1'b0;
    assign proc_15_start_FIFO_blk[2] = 1'b0;
    assign proc_15_TLF_FIFO_blk[2] = 1'b0;
    assign proc_15_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_15_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_15[2] = dl_detect_out ? proc_dep_vld_vec_15_reg[2] : (proc_15_data_FIFO_blk[2] | proc_15_data_PIPO_blk[2] | proc_15_start_FIFO_blk[2] | proc_15_TLF_FIFO_blk[2] | proc_15_input_sync_blk[2] | proc_15_output_sync_blk[2]);
    assign proc_15_data_FIFO_blk[3] = 1'b0;
    assign proc_15_data_PIPO_blk[3] = 1'b0;
    assign proc_15_start_FIFO_blk[3] = 1'b0;
    assign proc_15_TLF_FIFO_blk[3] = 1'b0;
    assign proc_15_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_15_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_15[3] = dl_detect_out ? proc_dep_vld_vec_15_reg[3] : (proc_15_data_FIFO_blk[3] | proc_15_data_PIPO_blk[3] | proc_15_start_FIFO_blk[3] | proc_15_TLF_FIFO_blk[3] | proc_15_input_sync_blk[3] | proc_15_output_sync_blk[3]);
    assign proc_15_data_FIFO_blk[4] = 1'b0;
    assign proc_15_data_PIPO_blk[4] = 1'b0;
    assign proc_15_start_FIFO_blk[4] = 1'b0;
    assign proc_15_TLF_FIFO_blk[4] = 1'b0;
    assign proc_15_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_15_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_15[4] = dl_detect_out ? proc_dep_vld_vec_15_reg[4] : (proc_15_data_FIFO_blk[4] | proc_15_data_PIPO_blk[4] | proc_15_start_FIFO_blk[4] | proc_15_TLF_FIFO_blk[4] | proc_15_input_sync_blk[4] | proc_15_output_sync_blk[4]);
    assign proc_15_data_FIFO_blk[5] = 1'b0;
    assign proc_15_data_PIPO_blk[5] = 1'b0;
    assign proc_15_start_FIFO_blk[5] = 1'b0;
    assign proc_15_TLF_FIFO_blk[5] = 1'b0;
    assign proc_15_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_15_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_15[5] = dl_detect_out ? proc_dep_vld_vec_15_reg[5] : (proc_15_data_FIFO_blk[5] | proc_15_data_PIPO_blk[5] | proc_15_start_FIFO_blk[5] | proc_15_TLF_FIFO_blk[5] | proc_15_input_sync_blk[5] | proc_15_output_sync_blk[5]);
    assign proc_15_data_FIFO_blk[6] = 1'b0;
    assign proc_15_data_PIPO_blk[6] = 1'b0;
    assign proc_15_start_FIFO_blk[6] = 1'b0;
    assign proc_15_TLF_FIFO_blk[6] = 1'b0;
    assign proc_15_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_15_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_15[6] = dl_detect_out ? proc_dep_vld_vec_15_reg[6] : (proc_15_data_FIFO_blk[6] | proc_15_data_PIPO_blk[6] | proc_15_start_FIFO_blk[6] | proc_15_TLF_FIFO_blk[6] | proc_15_input_sync_blk[6] | proc_15_output_sync_blk[6]);
    assign proc_15_data_FIFO_blk[7] = 1'b0;
    assign proc_15_data_PIPO_blk[7] = 1'b0;
    assign proc_15_start_FIFO_blk[7] = 1'b0;
    assign proc_15_TLF_FIFO_blk[7] = 1'b0;
    assign proc_15_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_15_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_15[7] = dl_detect_out ? proc_dep_vld_vec_15_reg[7] : (proc_15_data_FIFO_blk[7] | proc_15_data_PIPO_blk[7] | proc_15_start_FIFO_blk[7] | proc_15_TLF_FIFO_blk[7] | proc_15_input_sync_blk[7] | proc_15_output_sync_blk[7]);
    assign proc_15_data_FIFO_blk[8] = 1'b0;
    assign proc_15_data_PIPO_blk[8] = 1'b0;
    assign proc_15_start_FIFO_blk[8] = 1'b0;
    assign proc_15_TLF_FIFO_blk[8] = 1'b0;
    assign proc_15_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_15_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_15[8] = dl_detect_out ? proc_dep_vld_vec_15_reg[8] : (proc_15_data_FIFO_blk[8] | proc_15_data_PIPO_blk[8] | proc_15_start_FIFO_blk[8] | proc_15_TLF_FIFO_blk[8] | proc_15_input_sync_blk[8] | proc_15_output_sync_blk[8]);
    assign proc_15_data_FIFO_blk[9] = 1'b0;
    assign proc_15_data_PIPO_blk[9] = 1'b0;
    assign proc_15_start_FIFO_blk[9] = 1'b0;
    assign proc_15_TLF_FIFO_blk[9] = 1'b0;
    assign proc_15_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_15_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_15[9] = dl_detect_out ? proc_dep_vld_vec_15_reg[9] : (proc_15_data_FIFO_blk[9] | proc_15_data_PIPO_blk[9] | proc_15_start_FIFO_blk[9] | proc_15_TLF_FIFO_blk[9] | proc_15_input_sync_blk[9] | proc_15_output_sync_blk[9]);
    assign proc_15_data_FIFO_blk[10] = 1'b0;
    assign proc_15_data_PIPO_blk[10] = 1'b0;
    assign proc_15_start_FIFO_blk[10] = 1'b0;
    assign proc_15_TLF_FIFO_blk[10] = 1'b0;
    assign proc_15_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_15_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_15[10] = dl_detect_out ? proc_dep_vld_vec_15_reg[10] : (proc_15_data_FIFO_blk[10] | proc_15_data_PIPO_blk[10] | proc_15_start_FIFO_blk[10] | proc_15_TLF_FIFO_blk[10] | proc_15_input_sync_blk[10] | proc_15_output_sync_blk[10]);
    assign proc_15_data_FIFO_blk[11] = 1'b0;
    assign proc_15_data_PIPO_blk[11] = 1'b0;
    assign proc_15_start_FIFO_blk[11] = 1'b0;
    assign proc_15_TLF_FIFO_blk[11] = 1'b0;
    assign proc_15_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_15_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_15[11] = dl_detect_out ? proc_dep_vld_vec_15_reg[11] : (proc_15_data_FIFO_blk[11] | proc_15_data_PIPO_blk[11] | proc_15_start_FIFO_blk[11] | proc_15_TLF_FIFO_blk[11] | proc_15_input_sync_blk[11] | proc_15_output_sync_blk[11]);
    assign proc_15_data_FIFO_blk[12] = 1'b0;
    assign proc_15_data_PIPO_blk[12] = 1'b0;
    assign proc_15_start_FIFO_blk[12] = 1'b0;
    assign proc_15_TLF_FIFO_blk[12] = 1'b0;
    assign proc_15_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_15_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_15[12] = dl_detect_out ? proc_dep_vld_vec_15_reg[12] : (proc_15_data_FIFO_blk[12] | proc_15_data_PIPO_blk[12] | proc_15_start_FIFO_blk[12] | proc_15_TLF_FIFO_blk[12] | proc_15_input_sync_blk[12] | proc_15_output_sync_blk[12]);
    assign proc_15_data_FIFO_blk[13] = 1'b0;
    assign proc_15_data_PIPO_blk[13] = 1'b0;
    assign proc_15_start_FIFO_blk[13] = 1'b0;
    assign proc_15_TLF_FIFO_blk[13] = 1'b0;
    assign proc_15_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_15_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_15[13] = dl_detect_out ? proc_dep_vld_vec_15_reg[13] : (proc_15_data_FIFO_blk[13] | proc_15_data_PIPO_blk[13] | proc_15_start_FIFO_blk[13] | proc_15_TLF_FIFO_blk[13] | proc_15_input_sync_blk[13] | proc_15_output_sync_blk[13]);
    assign proc_15_data_FIFO_blk[14] = 1'b0;
    assign proc_15_data_PIPO_blk[14] = 1'b0;
    assign proc_15_start_FIFO_blk[14] = 1'b0;
    assign proc_15_TLF_FIFO_blk[14] = 1'b0;
    assign proc_15_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_15_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_15[14] = dl_detect_out ? proc_dep_vld_vec_15_reg[14] : (proc_15_data_FIFO_blk[14] | proc_15_data_PIPO_blk[14] | proc_15_start_FIFO_blk[14] | proc_15_TLF_FIFO_blk[14] | proc_15_input_sync_blk[14] | proc_15_output_sync_blk[14]);
    assign proc_15_data_FIFO_blk[15] = 1'b0;
    assign proc_15_data_PIPO_blk[15] = 1'b0;
    assign proc_15_start_FIFO_blk[15] = 1'b0;
    assign proc_15_TLF_FIFO_blk[15] = 1'b0;
    assign proc_15_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_15_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_15[15] = dl_detect_out ? proc_dep_vld_vec_15_reg[15] : (proc_15_data_FIFO_blk[15] | proc_15_data_PIPO_blk[15] | proc_15_start_FIFO_blk[15] | proc_15_TLF_FIFO_blk[15] | proc_15_input_sync_blk[15] | proc_15_output_sync_blk[15]);
    assign proc_15_data_FIFO_blk[16] = 1'b0;
    assign proc_15_data_PIPO_blk[16] = 1'b0;
    assign proc_15_start_FIFO_blk[16] = 1'b0;
    assign proc_15_TLF_FIFO_blk[16] = 1'b0;
    assign proc_15_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_15_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_15[16] = dl_detect_out ? proc_dep_vld_vec_15_reg[16] : (proc_15_data_FIFO_blk[16] | proc_15_data_PIPO_blk[16] | proc_15_start_FIFO_blk[16] | proc_15_TLF_FIFO_blk[16] | proc_15_input_sync_blk[16] | proc_15_output_sync_blk[16]);
    assign proc_15_data_FIFO_blk[17] = 1'b0;
    assign proc_15_data_PIPO_blk[17] = 1'b0;
    assign proc_15_start_FIFO_blk[17] = 1'b0;
    assign proc_15_TLF_FIFO_blk[17] = 1'b0;
    assign proc_15_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_15_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_15[17] = dl_detect_out ? proc_dep_vld_vec_15_reg[17] : (proc_15_data_FIFO_blk[17] | proc_15_data_PIPO_blk[17] | proc_15_start_FIFO_blk[17] | proc_15_TLF_FIFO_blk[17] | proc_15_input_sync_blk[17] | proc_15_output_sync_blk[17]);
    assign proc_15_data_FIFO_blk[18] = 1'b0;
    assign proc_15_data_PIPO_blk[18] = 1'b0;
    assign proc_15_start_FIFO_blk[18] = 1'b0;
    assign proc_15_TLF_FIFO_blk[18] = 1'b0;
    assign proc_15_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_15_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_15[18] = dl_detect_out ? proc_dep_vld_vec_15_reg[18] : (proc_15_data_FIFO_blk[18] | proc_15_data_PIPO_blk[18] | proc_15_start_FIFO_blk[18] | proc_15_TLF_FIFO_blk[18] | proc_15_input_sync_blk[18] | proc_15_output_sync_blk[18]);
    assign proc_15_data_FIFO_blk[19] = 1'b0;
    assign proc_15_data_PIPO_blk[19] = 1'b0;
    assign proc_15_start_FIFO_blk[19] = 1'b0;
    assign proc_15_TLF_FIFO_blk[19] = 1'b0;
    assign proc_15_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_15_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_15[19] = dl_detect_out ? proc_dep_vld_vec_15_reg[19] : (proc_15_data_FIFO_blk[19] | proc_15_data_PIPO_blk[19] | proc_15_start_FIFO_blk[19] | proc_15_TLF_FIFO_blk[19] | proc_15_input_sync_blk[19] | proc_15_output_sync_blk[19]);
    assign proc_15_data_FIFO_blk[20] = 1'b0;
    assign proc_15_data_PIPO_blk[20] = 1'b0;
    assign proc_15_start_FIFO_blk[20] = 1'b0;
    assign proc_15_TLF_FIFO_blk[20] = 1'b0;
    assign proc_15_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_15_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_15[20] = dl_detect_out ? proc_dep_vld_vec_15_reg[20] : (proc_15_data_FIFO_blk[20] | proc_15_data_PIPO_blk[20] | proc_15_start_FIFO_blk[20] | proc_15_TLF_FIFO_blk[20] | proc_15_input_sync_blk[20] | proc_15_output_sync_blk[20]);
    assign proc_15_data_FIFO_blk[21] = 1'b0;
    assign proc_15_data_PIPO_blk[21] = 1'b0;
    assign proc_15_start_FIFO_blk[21] = 1'b0;
    assign proc_15_TLF_FIFO_blk[21] = 1'b0;
    assign proc_15_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_15_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_15[21] = dl_detect_out ? proc_dep_vld_vec_15_reg[21] : (proc_15_data_FIFO_blk[21] | proc_15_data_PIPO_blk[21] | proc_15_start_FIFO_blk[21] | proc_15_TLF_FIFO_blk[21] | proc_15_input_sync_blk[21] | proc_15_output_sync_blk[21]);
    assign proc_15_data_FIFO_blk[22] = 1'b0;
    assign proc_15_data_PIPO_blk[22] = 1'b0;
    assign proc_15_start_FIFO_blk[22] = 1'b0;
    assign proc_15_TLF_FIFO_blk[22] = 1'b0;
    assign proc_15_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_15_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_15[22] = dl_detect_out ? proc_dep_vld_vec_15_reg[22] : (proc_15_data_FIFO_blk[22] | proc_15_data_PIPO_blk[22] | proc_15_start_FIFO_blk[22] | proc_15_TLF_FIFO_blk[22] | proc_15_input_sync_blk[22] | proc_15_output_sync_blk[22]);
    assign proc_15_data_FIFO_blk[23] = 1'b0;
    assign proc_15_data_PIPO_blk[23] = 1'b0;
    assign proc_15_start_FIFO_blk[23] = 1'b0;
    assign proc_15_TLF_FIFO_blk[23] = 1'b0;
    assign proc_15_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_15_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_15[23] = dl_detect_out ? proc_dep_vld_vec_15_reg[23] : (proc_15_data_FIFO_blk[23] | proc_15_data_PIPO_blk[23] | proc_15_start_FIFO_blk[23] | proc_15_TLF_FIFO_blk[23] | proc_15_input_sync_blk[23] | proc_15_output_sync_blk[23]);
    assign proc_15_data_FIFO_blk[24] = 1'b0;
    assign proc_15_data_PIPO_blk[24] = 1'b0;
    assign proc_15_start_FIFO_blk[24] = 1'b0;
    assign proc_15_TLF_FIFO_blk[24] = 1'b0;
    assign proc_15_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_15_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_15[24] = dl_detect_out ? proc_dep_vld_vec_15_reg[24] : (proc_15_data_FIFO_blk[24] | proc_15_data_PIPO_blk[24] | proc_15_start_FIFO_blk[24] | proc_15_TLF_FIFO_blk[24] | proc_15_input_sync_blk[24] | proc_15_output_sync_blk[24]);
    assign proc_15_data_FIFO_blk[25] = 1'b0;
    assign proc_15_data_PIPO_blk[25] = 1'b0;
    assign proc_15_start_FIFO_blk[25] = 1'b0;
    assign proc_15_TLF_FIFO_blk[25] = 1'b0;
    assign proc_15_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_15_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_15[25] = dl_detect_out ? proc_dep_vld_vec_15_reg[25] : (proc_15_data_FIFO_blk[25] | proc_15_data_PIPO_blk[25] | proc_15_start_FIFO_blk[25] | proc_15_TLF_FIFO_blk[25] | proc_15_input_sync_blk[25] | proc_15_output_sync_blk[25]);
    assign proc_15_data_FIFO_blk[26] = 1'b0;
    assign proc_15_data_PIPO_blk[26] = 1'b0;
    assign proc_15_start_FIFO_blk[26] = 1'b0;
    assign proc_15_TLF_FIFO_blk[26] = 1'b0;
    assign proc_15_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_15_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_15[26] = dl_detect_out ? proc_dep_vld_vec_15_reg[26] : (proc_15_data_FIFO_blk[26] | proc_15_data_PIPO_blk[26] | proc_15_start_FIFO_blk[26] | proc_15_TLF_FIFO_blk[26] | proc_15_input_sync_blk[26] | proc_15_output_sync_blk[26]);
    assign proc_15_data_FIFO_blk[27] = 1'b0;
    assign proc_15_data_PIPO_blk[27] = 1'b0;
    assign proc_15_start_FIFO_blk[27] = 1'b0;
    assign proc_15_TLF_FIFO_blk[27] = 1'b0;
    assign proc_15_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_15_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_15[27] = dl_detect_out ? proc_dep_vld_vec_15_reg[27] : (proc_15_data_FIFO_blk[27] | proc_15_data_PIPO_blk[27] | proc_15_start_FIFO_blk[27] | proc_15_TLF_FIFO_blk[27] | proc_15_input_sync_blk[27] | proc_15_output_sync_blk[27]);
    assign proc_15_data_FIFO_blk[28] = 1'b0;
    assign proc_15_data_PIPO_blk[28] = 1'b0;
    assign proc_15_start_FIFO_blk[28] = 1'b0;
    assign proc_15_TLF_FIFO_blk[28] = 1'b0;
    assign proc_15_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_15_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_15[28] = dl_detect_out ? proc_dep_vld_vec_15_reg[28] : (proc_15_data_FIFO_blk[28] | proc_15_data_PIPO_blk[28] | proc_15_start_FIFO_blk[28] | proc_15_TLF_FIFO_blk[28] | proc_15_input_sync_blk[28] | proc_15_output_sync_blk[28]);
    assign proc_15_data_FIFO_blk[29] = 1'b0;
    assign proc_15_data_PIPO_blk[29] = 1'b0;
    assign proc_15_start_FIFO_blk[29] = 1'b0;
    assign proc_15_TLF_FIFO_blk[29] = 1'b0;
    assign proc_15_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_15_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_15[29] = dl_detect_out ? proc_dep_vld_vec_15_reg[29] : (proc_15_data_FIFO_blk[29] | proc_15_data_PIPO_blk[29] | proc_15_start_FIFO_blk[29] | proc_15_TLF_FIFO_blk[29] | proc_15_input_sync_blk[29] | proc_15_output_sync_blk[29]);
    assign proc_15_data_FIFO_blk[30] = 1'b0;
    assign proc_15_data_PIPO_blk[30] = 1'b0;
    assign proc_15_start_FIFO_blk[30] = 1'b0;
    assign proc_15_TLF_FIFO_blk[30] = 1'b0;
    assign proc_15_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_15_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_15[30] = dl_detect_out ? proc_dep_vld_vec_15_reg[30] : (proc_15_data_FIFO_blk[30] | proc_15_data_PIPO_blk[30] | proc_15_start_FIFO_blk[30] | proc_15_TLF_FIFO_blk[30] | proc_15_input_sync_blk[30] | proc_15_output_sync_blk[30]);
    assign proc_15_data_FIFO_blk[31] = 1'b0;
    assign proc_15_data_PIPO_blk[31] = 1'b0;
    assign proc_15_start_FIFO_blk[31] = 1'b0;
    assign proc_15_TLF_FIFO_blk[31] = 1'b0;
    assign proc_15_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_15_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_15[31] = dl_detect_out ? proc_dep_vld_vec_15_reg[31] : (proc_15_data_FIFO_blk[31] | proc_15_data_PIPO_blk[31] | proc_15_start_FIFO_blk[31] | proc_15_TLF_FIFO_blk[31] | proc_15_input_sync_blk[31] | proc_15_output_sync_blk[31]);
    assign proc_15_data_FIFO_blk[32] = 1'b0;
    assign proc_15_data_PIPO_blk[32] = 1'b0;
    assign proc_15_start_FIFO_blk[32] = 1'b0;
    assign proc_15_TLF_FIFO_blk[32] = 1'b0;
    assign proc_15_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_10_U0_ap_ready & ProcessingElement_10_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_15_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_15[32] = dl_detect_out ? proc_dep_vld_vec_15_reg[32] : (proc_15_data_FIFO_blk[32] | proc_15_data_PIPO_blk[32] | proc_15_start_FIFO_blk[32] | proc_15_TLF_FIFO_blk[32] | proc_15_input_sync_blk[32] | proc_15_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_15_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_15_reg <= proc_dep_vld_vec_15;
        end
    end
    assign in_chan_dep_vld_vec_15[0] = dep_chan_vld_0_15;
    assign in_chan_dep_data_vec_15[39 : 0] = dep_chan_data_0_15;
    assign token_in_vec_15[0] = token_0_15;
    assign in_chan_dep_vld_vec_15[1] = dep_chan_vld_1_15;
    assign in_chan_dep_data_vec_15[79 : 40] = dep_chan_data_1_15;
    assign token_in_vec_15[1] = token_1_15;
    assign in_chan_dep_vld_vec_15[2] = dep_chan_vld_3_15;
    assign in_chan_dep_data_vec_15[119 : 80] = dep_chan_data_3_15;
    assign token_in_vec_15[2] = token_3_15;
    assign in_chan_dep_vld_vec_15[3] = dep_chan_vld_6_15;
    assign in_chan_dep_data_vec_15[159 : 120] = dep_chan_data_6_15;
    assign token_in_vec_15[3] = token_6_15;
    assign in_chan_dep_vld_vec_15[4] = dep_chan_vld_7_15;
    assign in_chan_dep_data_vec_15[199 : 160] = dep_chan_data_7_15;
    assign token_in_vec_15[4] = token_7_15;
    assign in_chan_dep_vld_vec_15[5] = dep_chan_vld_8_15;
    assign in_chan_dep_data_vec_15[239 : 200] = dep_chan_data_8_15;
    assign token_in_vec_15[5] = token_8_15;
    assign in_chan_dep_vld_vec_15[6] = dep_chan_vld_9_15;
    assign in_chan_dep_data_vec_15[279 : 240] = dep_chan_data_9_15;
    assign token_in_vec_15[6] = token_9_15;
    assign in_chan_dep_vld_vec_15[7] = dep_chan_vld_10_15;
    assign in_chan_dep_data_vec_15[319 : 280] = dep_chan_data_10_15;
    assign token_in_vec_15[7] = token_10_15;
    assign in_chan_dep_vld_vec_15[8] = dep_chan_vld_11_15;
    assign in_chan_dep_data_vec_15[359 : 320] = dep_chan_data_11_15;
    assign token_in_vec_15[8] = token_11_15;
    assign in_chan_dep_vld_vec_15[9] = dep_chan_vld_12_15;
    assign in_chan_dep_data_vec_15[399 : 360] = dep_chan_data_12_15;
    assign token_in_vec_15[9] = token_12_15;
    assign in_chan_dep_vld_vec_15[10] = dep_chan_vld_13_15;
    assign in_chan_dep_data_vec_15[439 : 400] = dep_chan_data_13_15;
    assign token_in_vec_15[10] = token_13_15;
    assign in_chan_dep_vld_vec_15[11] = dep_chan_vld_14_15;
    assign in_chan_dep_data_vec_15[479 : 440] = dep_chan_data_14_15;
    assign token_in_vec_15[11] = token_14_15;
    assign in_chan_dep_vld_vec_15[12] = dep_chan_vld_16_15;
    assign in_chan_dep_data_vec_15[519 : 480] = dep_chan_data_16_15;
    assign token_in_vec_15[12] = token_16_15;
    assign in_chan_dep_vld_vec_15[13] = dep_chan_vld_17_15;
    assign in_chan_dep_data_vec_15[559 : 520] = dep_chan_data_17_15;
    assign token_in_vec_15[13] = token_17_15;
    assign in_chan_dep_vld_vec_15[14] = dep_chan_vld_18_15;
    assign in_chan_dep_data_vec_15[599 : 560] = dep_chan_data_18_15;
    assign token_in_vec_15[14] = token_18_15;
    assign in_chan_dep_vld_vec_15[15] = dep_chan_vld_19_15;
    assign in_chan_dep_data_vec_15[639 : 600] = dep_chan_data_19_15;
    assign token_in_vec_15[15] = token_19_15;
    assign in_chan_dep_vld_vec_15[16] = dep_chan_vld_20_15;
    assign in_chan_dep_data_vec_15[679 : 640] = dep_chan_data_20_15;
    assign token_in_vec_15[16] = token_20_15;
    assign in_chan_dep_vld_vec_15[17] = dep_chan_vld_21_15;
    assign in_chan_dep_data_vec_15[719 : 680] = dep_chan_data_21_15;
    assign token_in_vec_15[17] = token_21_15;
    assign in_chan_dep_vld_vec_15[18] = dep_chan_vld_22_15;
    assign in_chan_dep_data_vec_15[759 : 720] = dep_chan_data_22_15;
    assign token_in_vec_15[18] = token_22_15;
    assign in_chan_dep_vld_vec_15[19] = dep_chan_vld_23_15;
    assign in_chan_dep_data_vec_15[799 : 760] = dep_chan_data_23_15;
    assign token_in_vec_15[19] = token_23_15;
    assign in_chan_dep_vld_vec_15[20] = dep_chan_vld_24_15;
    assign in_chan_dep_data_vec_15[839 : 800] = dep_chan_data_24_15;
    assign token_in_vec_15[20] = token_24_15;
    assign in_chan_dep_vld_vec_15[21] = dep_chan_vld_25_15;
    assign in_chan_dep_data_vec_15[879 : 840] = dep_chan_data_25_15;
    assign token_in_vec_15[21] = token_25_15;
    assign in_chan_dep_vld_vec_15[22] = dep_chan_vld_26_15;
    assign in_chan_dep_data_vec_15[919 : 880] = dep_chan_data_26_15;
    assign token_in_vec_15[22] = token_26_15;
    assign in_chan_dep_vld_vec_15[23] = dep_chan_vld_27_15;
    assign in_chan_dep_data_vec_15[959 : 920] = dep_chan_data_27_15;
    assign token_in_vec_15[23] = token_27_15;
    assign in_chan_dep_vld_vec_15[24] = dep_chan_vld_28_15;
    assign in_chan_dep_data_vec_15[999 : 960] = dep_chan_data_28_15;
    assign token_in_vec_15[24] = token_28_15;
    assign in_chan_dep_vld_vec_15[25] = dep_chan_vld_29_15;
    assign in_chan_dep_data_vec_15[1039 : 1000] = dep_chan_data_29_15;
    assign token_in_vec_15[25] = token_29_15;
    assign in_chan_dep_vld_vec_15[26] = dep_chan_vld_30_15;
    assign in_chan_dep_data_vec_15[1079 : 1040] = dep_chan_data_30_15;
    assign token_in_vec_15[26] = token_30_15;
    assign in_chan_dep_vld_vec_15[27] = dep_chan_vld_31_15;
    assign in_chan_dep_data_vec_15[1119 : 1080] = dep_chan_data_31_15;
    assign token_in_vec_15[27] = token_31_15;
    assign in_chan_dep_vld_vec_15[28] = dep_chan_vld_32_15;
    assign in_chan_dep_data_vec_15[1159 : 1120] = dep_chan_data_32_15;
    assign token_in_vec_15[28] = token_32_15;
    assign in_chan_dep_vld_vec_15[29] = dep_chan_vld_33_15;
    assign in_chan_dep_data_vec_15[1199 : 1160] = dep_chan_data_33_15;
    assign token_in_vec_15[29] = token_33_15;
    assign in_chan_dep_vld_vec_15[30] = dep_chan_vld_34_15;
    assign in_chan_dep_data_vec_15[1239 : 1200] = dep_chan_data_34_15;
    assign token_in_vec_15[30] = token_34_15;
    assign in_chan_dep_vld_vec_15[31] = dep_chan_vld_35_15;
    assign in_chan_dep_data_vec_15[1279 : 1240] = dep_chan_data_35_15;
    assign token_in_vec_15[31] = token_35_15;
    assign in_chan_dep_vld_vec_15[32] = dep_chan_vld_36_15;
    assign in_chan_dep_data_vec_15[1319 : 1280] = dep_chan_data_36_15;
    assign token_in_vec_15[32] = token_36_15;
    assign dep_chan_vld_15_14 = out_chan_dep_vld_vec_15[0];
    assign dep_chan_data_15_14 = out_chan_dep_data_15;
    assign token_15_14 = token_out_vec_15[0];
    assign dep_chan_vld_15_16 = out_chan_dep_vld_vec_15[1];
    assign dep_chan_data_15_16 = out_chan_dep_data_15;
    assign token_15_16 = token_out_vec_15[1];
    assign dep_chan_vld_15_0 = out_chan_dep_vld_vec_15[2];
    assign dep_chan_data_15_0 = out_chan_dep_data_15;
    assign token_15_0 = token_out_vec_15[2];
    assign dep_chan_vld_15_1 = out_chan_dep_vld_vec_15[3];
    assign dep_chan_data_15_1 = out_chan_dep_data_15;
    assign token_15_1 = token_out_vec_15[3];
    assign dep_chan_vld_15_3 = out_chan_dep_vld_vec_15[4];
    assign dep_chan_data_15_3 = out_chan_dep_data_15;
    assign token_15_3 = token_out_vec_15[4];
    assign dep_chan_vld_15_6 = out_chan_dep_vld_vec_15[5];
    assign dep_chan_data_15_6 = out_chan_dep_data_15;
    assign token_15_6 = token_out_vec_15[5];
    assign dep_chan_vld_15_7 = out_chan_dep_vld_vec_15[6];
    assign dep_chan_data_15_7 = out_chan_dep_data_15;
    assign token_15_7 = token_out_vec_15[6];
    assign dep_chan_vld_15_8 = out_chan_dep_vld_vec_15[7];
    assign dep_chan_data_15_8 = out_chan_dep_data_15;
    assign token_15_8 = token_out_vec_15[7];
    assign dep_chan_vld_15_9 = out_chan_dep_vld_vec_15[8];
    assign dep_chan_data_15_9 = out_chan_dep_data_15;
    assign token_15_9 = token_out_vec_15[8];
    assign dep_chan_vld_15_10 = out_chan_dep_vld_vec_15[9];
    assign dep_chan_data_15_10 = out_chan_dep_data_15;
    assign token_15_10 = token_out_vec_15[9];
    assign dep_chan_vld_15_11 = out_chan_dep_vld_vec_15[10];
    assign dep_chan_data_15_11 = out_chan_dep_data_15;
    assign token_15_11 = token_out_vec_15[10];
    assign dep_chan_vld_15_12 = out_chan_dep_vld_vec_15[11];
    assign dep_chan_data_15_12 = out_chan_dep_data_15;
    assign token_15_12 = token_out_vec_15[11];
    assign dep_chan_vld_15_13 = out_chan_dep_vld_vec_15[12];
    assign dep_chan_data_15_13 = out_chan_dep_data_15;
    assign token_15_13 = token_out_vec_15[12];
    assign dep_chan_vld_15_17 = out_chan_dep_vld_vec_15[13];
    assign dep_chan_data_15_17 = out_chan_dep_data_15;
    assign token_15_17 = token_out_vec_15[13];
    assign dep_chan_vld_15_18 = out_chan_dep_vld_vec_15[14];
    assign dep_chan_data_15_18 = out_chan_dep_data_15;
    assign token_15_18 = token_out_vec_15[14];
    assign dep_chan_vld_15_19 = out_chan_dep_vld_vec_15[15];
    assign dep_chan_data_15_19 = out_chan_dep_data_15;
    assign token_15_19 = token_out_vec_15[15];
    assign dep_chan_vld_15_20 = out_chan_dep_vld_vec_15[16];
    assign dep_chan_data_15_20 = out_chan_dep_data_15;
    assign token_15_20 = token_out_vec_15[16];
    assign dep_chan_vld_15_21 = out_chan_dep_vld_vec_15[17];
    assign dep_chan_data_15_21 = out_chan_dep_data_15;
    assign token_15_21 = token_out_vec_15[17];
    assign dep_chan_vld_15_22 = out_chan_dep_vld_vec_15[18];
    assign dep_chan_data_15_22 = out_chan_dep_data_15;
    assign token_15_22 = token_out_vec_15[18];
    assign dep_chan_vld_15_23 = out_chan_dep_vld_vec_15[19];
    assign dep_chan_data_15_23 = out_chan_dep_data_15;
    assign token_15_23 = token_out_vec_15[19];
    assign dep_chan_vld_15_24 = out_chan_dep_vld_vec_15[20];
    assign dep_chan_data_15_24 = out_chan_dep_data_15;
    assign token_15_24 = token_out_vec_15[20];
    assign dep_chan_vld_15_25 = out_chan_dep_vld_vec_15[21];
    assign dep_chan_data_15_25 = out_chan_dep_data_15;
    assign token_15_25 = token_out_vec_15[21];
    assign dep_chan_vld_15_26 = out_chan_dep_vld_vec_15[22];
    assign dep_chan_data_15_26 = out_chan_dep_data_15;
    assign token_15_26 = token_out_vec_15[22];
    assign dep_chan_vld_15_27 = out_chan_dep_vld_vec_15[23];
    assign dep_chan_data_15_27 = out_chan_dep_data_15;
    assign token_15_27 = token_out_vec_15[23];
    assign dep_chan_vld_15_28 = out_chan_dep_vld_vec_15[24];
    assign dep_chan_data_15_28 = out_chan_dep_data_15;
    assign token_15_28 = token_out_vec_15[24];
    assign dep_chan_vld_15_29 = out_chan_dep_vld_vec_15[25];
    assign dep_chan_data_15_29 = out_chan_dep_data_15;
    assign token_15_29 = token_out_vec_15[25];
    assign dep_chan_vld_15_30 = out_chan_dep_vld_vec_15[26];
    assign dep_chan_data_15_30 = out_chan_dep_data_15;
    assign token_15_30 = token_out_vec_15[26];
    assign dep_chan_vld_15_31 = out_chan_dep_vld_vec_15[27];
    assign dep_chan_data_15_31 = out_chan_dep_data_15;
    assign token_15_31 = token_out_vec_15[27];
    assign dep_chan_vld_15_32 = out_chan_dep_vld_vec_15[28];
    assign dep_chan_data_15_32 = out_chan_dep_data_15;
    assign token_15_32 = token_out_vec_15[28];
    assign dep_chan_vld_15_33 = out_chan_dep_vld_vec_15[29];
    assign dep_chan_data_15_33 = out_chan_dep_data_15;
    assign token_15_33 = token_out_vec_15[29];
    assign dep_chan_vld_15_34 = out_chan_dep_vld_vec_15[30];
    assign dep_chan_data_15_34 = out_chan_dep_data_15;
    assign token_15_34 = token_out_vec_15[30];
    assign dep_chan_vld_15_35 = out_chan_dep_vld_vec_15[31];
    assign dep_chan_data_15_35 = out_chan_dep_data_15;
    assign token_15_35 = token_out_vec_15[31];
    assign dep_chan_vld_15_36 = out_chan_dep_vld_vec_15[32];
    assign dep_chan_data_15_36 = out_chan_dep_data_15;
    assign token_15_36 = token_out_vec_15[32];

    // Process: ProcessingElement_11_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 16, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_16 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_16),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_16),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_16),
        .token_in_vec(token_in_vec_16),
        .dl_detect_in(dl_detect_out),
        .origin(origin[16]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_16),
        .out_chan_dep_data(out_chan_dep_data_16),
        .token_out_vec(token_out_vec_16),
        .dl_detect_out(dl_in_vec[16]));

    assign proc_16_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_10_blk_n) | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_10_blk_n) | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_WriteC_Flattened_fu_179.cPipes_10_blk_n);
    assign proc_16_data_PIPO_blk[0] = 1'b0;
    assign proc_16_start_FIFO_blk[0] = 1'b0;
    assign proc_16_TLF_FIFO_blk[0] = 1'b0;
    assign proc_16_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_16_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_16[0] = dl_detect_out ? proc_dep_vld_vec_16_reg[0] : (proc_16_data_FIFO_blk[0] | proc_16_data_PIPO_blk[0] | proc_16_start_FIFO_blk[0] | proc_16_TLF_FIFO_blk[0] | proc_16_input_sync_blk[0] | proc_16_output_sync_blk[0]);
    assign proc_16_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_11_blk_n) | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_11_blk_n) | (~ProcessingElement_11_U0.grp_ProcessingElement_11_Pipeline_WriteC_Flattened_fu_179.cPipes_11_blk_n);
    assign proc_16_data_PIPO_blk[1] = 1'b0;
    assign proc_16_start_FIFO_blk[1] = 1'b0;
    assign proc_16_TLF_FIFO_blk[1] = 1'b0;
    assign proc_16_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_16_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_16[1] = dl_detect_out ? proc_dep_vld_vec_16_reg[1] : (proc_16_data_FIFO_blk[1] | proc_16_data_PIPO_blk[1] | proc_16_start_FIFO_blk[1] | proc_16_TLF_FIFO_blk[1] | proc_16_input_sync_blk[1] | proc_16_output_sync_blk[1]);
    assign proc_16_data_FIFO_blk[2] = 1'b0;
    assign proc_16_data_PIPO_blk[2] = 1'b0;
    assign proc_16_start_FIFO_blk[2] = 1'b0;
    assign proc_16_TLF_FIFO_blk[2] = 1'b0;
    assign proc_16_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_16_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_16[2] = dl_detect_out ? proc_dep_vld_vec_16_reg[2] : (proc_16_data_FIFO_blk[2] | proc_16_data_PIPO_blk[2] | proc_16_start_FIFO_blk[2] | proc_16_TLF_FIFO_blk[2] | proc_16_input_sync_blk[2] | proc_16_output_sync_blk[2]);
    assign proc_16_data_FIFO_blk[3] = 1'b0;
    assign proc_16_data_PIPO_blk[3] = 1'b0;
    assign proc_16_start_FIFO_blk[3] = 1'b0;
    assign proc_16_TLF_FIFO_blk[3] = 1'b0;
    assign proc_16_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_16_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_16[3] = dl_detect_out ? proc_dep_vld_vec_16_reg[3] : (proc_16_data_FIFO_blk[3] | proc_16_data_PIPO_blk[3] | proc_16_start_FIFO_blk[3] | proc_16_TLF_FIFO_blk[3] | proc_16_input_sync_blk[3] | proc_16_output_sync_blk[3]);
    assign proc_16_data_FIFO_blk[4] = 1'b0;
    assign proc_16_data_PIPO_blk[4] = 1'b0;
    assign proc_16_start_FIFO_blk[4] = 1'b0;
    assign proc_16_TLF_FIFO_blk[4] = 1'b0;
    assign proc_16_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_16_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_16[4] = dl_detect_out ? proc_dep_vld_vec_16_reg[4] : (proc_16_data_FIFO_blk[4] | proc_16_data_PIPO_blk[4] | proc_16_start_FIFO_blk[4] | proc_16_TLF_FIFO_blk[4] | proc_16_input_sync_blk[4] | proc_16_output_sync_blk[4]);
    assign proc_16_data_FIFO_blk[5] = 1'b0;
    assign proc_16_data_PIPO_blk[5] = 1'b0;
    assign proc_16_start_FIFO_blk[5] = 1'b0;
    assign proc_16_TLF_FIFO_blk[5] = 1'b0;
    assign proc_16_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_16_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_16[5] = dl_detect_out ? proc_dep_vld_vec_16_reg[5] : (proc_16_data_FIFO_blk[5] | proc_16_data_PIPO_blk[5] | proc_16_start_FIFO_blk[5] | proc_16_TLF_FIFO_blk[5] | proc_16_input_sync_blk[5] | proc_16_output_sync_blk[5]);
    assign proc_16_data_FIFO_blk[6] = 1'b0;
    assign proc_16_data_PIPO_blk[6] = 1'b0;
    assign proc_16_start_FIFO_blk[6] = 1'b0;
    assign proc_16_TLF_FIFO_blk[6] = 1'b0;
    assign proc_16_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_16_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_16[6] = dl_detect_out ? proc_dep_vld_vec_16_reg[6] : (proc_16_data_FIFO_blk[6] | proc_16_data_PIPO_blk[6] | proc_16_start_FIFO_blk[6] | proc_16_TLF_FIFO_blk[6] | proc_16_input_sync_blk[6] | proc_16_output_sync_blk[6]);
    assign proc_16_data_FIFO_blk[7] = 1'b0;
    assign proc_16_data_PIPO_blk[7] = 1'b0;
    assign proc_16_start_FIFO_blk[7] = 1'b0;
    assign proc_16_TLF_FIFO_blk[7] = 1'b0;
    assign proc_16_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_16_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_16[7] = dl_detect_out ? proc_dep_vld_vec_16_reg[7] : (proc_16_data_FIFO_blk[7] | proc_16_data_PIPO_blk[7] | proc_16_start_FIFO_blk[7] | proc_16_TLF_FIFO_blk[7] | proc_16_input_sync_blk[7] | proc_16_output_sync_blk[7]);
    assign proc_16_data_FIFO_blk[8] = 1'b0;
    assign proc_16_data_PIPO_blk[8] = 1'b0;
    assign proc_16_start_FIFO_blk[8] = 1'b0;
    assign proc_16_TLF_FIFO_blk[8] = 1'b0;
    assign proc_16_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_16_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_16[8] = dl_detect_out ? proc_dep_vld_vec_16_reg[8] : (proc_16_data_FIFO_blk[8] | proc_16_data_PIPO_blk[8] | proc_16_start_FIFO_blk[8] | proc_16_TLF_FIFO_blk[8] | proc_16_input_sync_blk[8] | proc_16_output_sync_blk[8]);
    assign proc_16_data_FIFO_blk[9] = 1'b0;
    assign proc_16_data_PIPO_blk[9] = 1'b0;
    assign proc_16_start_FIFO_blk[9] = 1'b0;
    assign proc_16_TLF_FIFO_blk[9] = 1'b0;
    assign proc_16_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_16_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_16[9] = dl_detect_out ? proc_dep_vld_vec_16_reg[9] : (proc_16_data_FIFO_blk[9] | proc_16_data_PIPO_blk[9] | proc_16_start_FIFO_blk[9] | proc_16_TLF_FIFO_blk[9] | proc_16_input_sync_blk[9] | proc_16_output_sync_blk[9]);
    assign proc_16_data_FIFO_blk[10] = 1'b0;
    assign proc_16_data_PIPO_blk[10] = 1'b0;
    assign proc_16_start_FIFO_blk[10] = 1'b0;
    assign proc_16_TLF_FIFO_blk[10] = 1'b0;
    assign proc_16_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_16_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_16[10] = dl_detect_out ? proc_dep_vld_vec_16_reg[10] : (proc_16_data_FIFO_blk[10] | proc_16_data_PIPO_blk[10] | proc_16_start_FIFO_blk[10] | proc_16_TLF_FIFO_blk[10] | proc_16_input_sync_blk[10] | proc_16_output_sync_blk[10]);
    assign proc_16_data_FIFO_blk[11] = 1'b0;
    assign proc_16_data_PIPO_blk[11] = 1'b0;
    assign proc_16_start_FIFO_blk[11] = 1'b0;
    assign proc_16_TLF_FIFO_blk[11] = 1'b0;
    assign proc_16_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_16_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_16[11] = dl_detect_out ? proc_dep_vld_vec_16_reg[11] : (proc_16_data_FIFO_blk[11] | proc_16_data_PIPO_blk[11] | proc_16_start_FIFO_blk[11] | proc_16_TLF_FIFO_blk[11] | proc_16_input_sync_blk[11] | proc_16_output_sync_blk[11]);
    assign proc_16_data_FIFO_blk[12] = 1'b0;
    assign proc_16_data_PIPO_blk[12] = 1'b0;
    assign proc_16_start_FIFO_blk[12] = 1'b0;
    assign proc_16_TLF_FIFO_blk[12] = 1'b0;
    assign proc_16_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_16_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_16[12] = dl_detect_out ? proc_dep_vld_vec_16_reg[12] : (proc_16_data_FIFO_blk[12] | proc_16_data_PIPO_blk[12] | proc_16_start_FIFO_blk[12] | proc_16_TLF_FIFO_blk[12] | proc_16_input_sync_blk[12] | proc_16_output_sync_blk[12]);
    assign proc_16_data_FIFO_blk[13] = 1'b0;
    assign proc_16_data_PIPO_blk[13] = 1'b0;
    assign proc_16_start_FIFO_blk[13] = 1'b0;
    assign proc_16_TLF_FIFO_blk[13] = 1'b0;
    assign proc_16_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_16_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_16[13] = dl_detect_out ? proc_dep_vld_vec_16_reg[13] : (proc_16_data_FIFO_blk[13] | proc_16_data_PIPO_blk[13] | proc_16_start_FIFO_blk[13] | proc_16_TLF_FIFO_blk[13] | proc_16_input_sync_blk[13] | proc_16_output_sync_blk[13]);
    assign proc_16_data_FIFO_blk[14] = 1'b0;
    assign proc_16_data_PIPO_blk[14] = 1'b0;
    assign proc_16_start_FIFO_blk[14] = 1'b0;
    assign proc_16_TLF_FIFO_blk[14] = 1'b0;
    assign proc_16_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_16_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_16[14] = dl_detect_out ? proc_dep_vld_vec_16_reg[14] : (proc_16_data_FIFO_blk[14] | proc_16_data_PIPO_blk[14] | proc_16_start_FIFO_blk[14] | proc_16_TLF_FIFO_blk[14] | proc_16_input_sync_blk[14] | proc_16_output_sync_blk[14]);
    assign proc_16_data_FIFO_blk[15] = 1'b0;
    assign proc_16_data_PIPO_blk[15] = 1'b0;
    assign proc_16_start_FIFO_blk[15] = 1'b0;
    assign proc_16_TLF_FIFO_blk[15] = 1'b0;
    assign proc_16_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_16_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_16[15] = dl_detect_out ? proc_dep_vld_vec_16_reg[15] : (proc_16_data_FIFO_blk[15] | proc_16_data_PIPO_blk[15] | proc_16_start_FIFO_blk[15] | proc_16_TLF_FIFO_blk[15] | proc_16_input_sync_blk[15] | proc_16_output_sync_blk[15]);
    assign proc_16_data_FIFO_blk[16] = 1'b0;
    assign proc_16_data_PIPO_blk[16] = 1'b0;
    assign proc_16_start_FIFO_blk[16] = 1'b0;
    assign proc_16_TLF_FIFO_blk[16] = 1'b0;
    assign proc_16_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_16_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_16[16] = dl_detect_out ? proc_dep_vld_vec_16_reg[16] : (proc_16_data_FIFO_blk[16] | proc_16_data_PIPO_blk[16] | proc_16_start_FIFO_blk[16] | proc_16_TLF_FIFO_blk[16] | proc_16_input_sync_blk[16] | proc_16_output_sync_blk[16]);
    assign proc_16_data_FIFO_blk[17] = 1'b0;
    assign proc_16_data_PIPO_blk[17] = 1'b0;
    assign proc_16_start_FIFO_blk[17] = 1'b0;
    assign proc_16_TLF_FIFO_blk[17] = 1'b0;
    assign proc_16_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_16_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_16[17] = dl_detect_out ? proc_dep_vld_vec_16_reg[17] : (proc_16_data_FIFO_blk[17] | proc_16_data_PIPO_blk[17] | proc_16_start_FIFO_blk[17] | proc_16_TLF_FIFO_blk[17] | proc_16_input_sync_blk[17] | proc_16_output_sync_blk[17]);
    assign proc_16_data_FIFO_blk[18] = 1'b0;
    assign proc_16_data_PIPO_blk[18] = 1'b0;
    assign proc_16_start_FIFO_blk[18] = 1'b0;
    assign proc_16_TLF_FIFO_blk[18] = 1'b0;
    assign proc_16_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_16_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_16[18] = dl_detect_out ? proc_dep_vld_vec_16_reg[18] : (proc_16_data_FIFO_blk[18] | proc_16_data_PIPO_blk[18] | proc_16_start_FIFO_blk[18] | proc_16_TLF_FIFO_blk[18] | proc_16_input_sync_blk[18] | proc_16_output_sync_blk[18]);
    assign proc_16_data_FIFO_blk[19] = 1'b0;
    assign proc_16_data_PIPO_blk[19] = 1'b0;
    assign proc_16_start_FIFO_blk[19] = 1'b0;
    assign proc_16_TLF_FIFO_blk[19] = 1'b0;
    assign proc_16_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_16_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_16[19] = dl_detect_out ? proc_dep_vld_vec_16_reg[19] : (proc_16_data_FIFO_blk[19] | proc_16_data_PIPO_blk[19] | proc_16_start_FIFO_blk[19] | proc_16_TLF_FIFO_blk[19] | proc_16_input_sync_blk[19] | proc_16_output_sync_blk[19]);
    assign proc_16_data_FIFO_blk[20] = 1'b0;
    assign proc_16_data_PIPO_blk[20] = 1'b0;
    assign proc_16_start_FIFO_blk[20] = 1'b0;
    assign proc_16_TLF_FIFO_blk[20] = 1'b0;
    assign proc_16_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_16_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_16[20] = dl_detect_out ? proc_dep_vld_vec_16_reg[20] : (proc_16_data_FIFO_blk[20] | proc_16_data_PIPO_blk[20] | proc_16_start_FIFO_blk[20] | proc_16_TLF_FIFO_blk[20] | proc_16_input_sync_blk[20] | proc_16_output_sync_blk[20]);
    assign proc_16_data_FIFO_blk[21] = 1'b0;
    assign proc_16_data_PIPO_blk[21] = 1'b0;
    assign proc_16_start_FIFO_blk[21] = 1'b0;
    assign proc_16_TLF_FIFO_blk[21] = 1'b0;
    assign proc_16_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_16_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_16[21] = dl_detect_out ? proc_dep_vld_vec_16_reg[21] : (proc_16_data_FIFO_blk[21] | proc_16_data_PIPO_blk[21] | proc_16_start_FIFO_blk[21] | proc_16_TLF_FIFO_blk[21] | proc_16_input_sync_blk[21] | proc_16_output_sync_blk[21]);
    assign proc_16_data_FIFO_blk[22] = 1'b0;
    assign proc_16_data_PIPO_blk[22] = 1'b0;
    assign proc_16_start_FIFO_blk[22] = 1'b0;
    assign proc_16_TLF_FIFO_blk[22] = 1'b0;
    assign proc_16_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_16_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_16[22] = dl_detect_out ? proc_dep_vld_vec_16_reg[22] : (proc_16_data_FIFO_blk[22] | proc_16_data_PIPO_blk[22] | proc_16_start_FIFO_blk[22] | proc_16_TLF_FIFO_blk[22] | proc_16_input_sync_blk[22] | proc_16_output_sync_blk[22]);
    assign proc_16_data_FIFO_blk[23] = 1'b0;
    assign proc_16_data_PIPO_blk[23] = 1'b0;
    assign proc_16_start_FIFO_blk[23] = 1'b0;
    assign proc_16_TLF_FIFO_blk[23] = 1'b0;
    assign proc_16_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_16_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_16[23] = dl_detect_out ? proc_dep_vld_vec_16_reg[23] : (proc_16_data_FIFO_blk[23] | proc_16_data_PIPO_blk[23] | proc_16_start_FIFO_blk[23] | proc_16_TLF_FIFO_blk[23] | proc_16_input_sync_blk[23] | proc_16_output_sync_blk[23]);
    assign proc_16_data_FIFO_blk[24] = 1'b0;
    assign proc_16_data_PIPO_blk[24] = 1'b0;
    assign proc_16_start_FIFO_blk[24] = 1'b0;
    assign proc_16_TLF_FIFO_blk[24] = 1'b0;
    assign proc_16_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_16_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_16[24] = dl_detect_out ? proc_dep_vld_vec_16_reg[24] : (proc_16_data_FIFO_blk[24] | proc_16_data_PIPO_blk[24] | proc_16_start_FIFO_blk[24] | proc_16_TLF_FIFO_blk[24] | proc_16_input_sync_blk[24] | proc_16_output_sync_blk[24]);
    assign proc_16_data_FIFO_blk[25] = 1'b0;
    assign proc_16_data_PIPO_blk[25] = 1'b0;
    assign proc_16_start_FIFO_blk[25] = 1'b0;
    assign proc_16_TLF_FIFO_blk[25] = 1'b0;
    assign proc_16_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_16_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_16[25] = dl_detect_out ? proc_dep_vld_vec_16_reg[25] : (proc_16_data_FIFO_blk[25] | proc_16_data_PIPO_blk[25] | proc_16_start_FIFO_blk[25] | proc_16_TLF_FIFO_blk[25] | proc_16_input_sync_blk[25] | proc_16_output_sync_blk[25]);
    assign proc_16_data_FIFO_blk[26] = 1'b0;
    assign proc_16_data_PIPO_blk[26] = 1'b0;
    assign proc_16_start_FIFO_blk[26] = 1'b0;
    assign proc_16_TLF_FIFO_blk[26] = 1'b0;
    assign proc_16_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_16_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_16[26] = dl_detect_out ? proc_dep_vld_vec_16_reg[26] : (proc_16_data_FIFO_blk[26] | proc_16_data_PIPO_blk[26] | proc_16_start_FIFO_blk[26] | proc_16_TLF_FIFO_blk[26] | proc_16_input_sync_blk[26] | proc_16_output_sync_blk[26]);
    assign proc_16_data_FIFO_blk[27] = 1'b0;
    assign proc_16_data_PIPO_blk[27] = 1'b0;
    assign proc_16_start_FIFO_blk[27] = 1'b0;
    assign proc_16_TLF_FIFO_blk[27] = 1'b0;
    assign proc_16_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_16_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_16[27] = dl_detect_out ? proc_dep_vld_vec_16_reg[27] : (proc_16_data_FIFO_blk[27] | proc_16_data_PIPO_blk[27] | proc_16_start_FIFO_blk[27] | proc_16_TLF_FIFO_blk[27] | proc_16_input_sync_blk[27] | proc_16_output_sync_blk[27]);
    assign proc_16_data_FIFO_blk[28] = 1'b0;
    assign proc_16_data_PIPO_blk[28] = 1'b0;
    assign proc_16_start_FIFO_blk[28] = 1'b0;
    assign proc_16_TLF_FIFO_blk[28] = 1'b0;
    assign proc_16_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_16_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_16[28] = dl_detect_out ? proc_dep_vld_vec_16_reg[28] : (proc_16_data_FIFO_blk[28] | proc_16_data_PIPO_blk[28] | proc_16_start_FIFO_blk[28] | proc_16_TLF_FIFO_blk[28] | proc_16_input_sync_blk[28] | proc_16_output_sync_blk[28]);
    assign proc_16_data_FIFO_blk[29] = 1'b0;
    assign proc_16_data_PIPO_blk[29] = 1'b0;
    assign proc_16_start_FIFO_blk[29] = 1'b0;
    assign proc_16_TLF_FIFO_blk[29] = 1'b0;
    assign proc_16_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_16_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_16[29] = dl_detect_out ? proc_dep_vld_vec_16_reg[29] : (proc_16_data_FIFO_blk[29] | proc_16_data_PIPO_blk[29] | proc_16_start_FIFO_blk[29] | proc_16_TLF_FIFO_blk[29] | proc_16_input_sync_blk[29] | proc_16_output_sync_blk[29]);
    assign proc_16_data_FIFO_blk[30] = 1'b0;
    assign proc_16_data_PIPO_blk[30] = 1'b0;
    assign proc_16_start_FIFO_blk[30] = 1'b0;
    assign proc_16_TLF_FIFO_blk[30] = 1'b0;
    assign proc_16_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_16_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_16[30] = dl_detect_out ? proc_dep_vld_vec_16_reg[30] : (proc_16_data_FIFO_blk[30] | proc_16_data_PIPO_blk[30] | proc_16_start_FIFO_blk[30] | proc_16_TLF_FIFO_blk[30] | proc_16_input_sync_blk[30] | proc_16_output_sync_blk[30]);
    assign proc_16_data_FIFO_blk[31] = 1'b0;
    assign proc_16_data_PIPO_blk[31] = 1'b0;
    assign proc_16_start_FIFO_blk[31] = 1'b0;
    assign proc_16_TLF_FIFO_blk[31] = 1'b0;
    assign proc_16_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_16_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_16[31] = dl_detect_out ? proc_dep_vld_vec_16_reg[31] : (proc_16_data_FIFO_blk[31] | proc_16_data_PIPO_blk[31] | proc_16_start_FIFO_blk[31] | proc_16_TLF_FIFO_blk[31] | proc_16_input_sync_blk[31] | proc_16_output_sync_blk[31]);
    assign proc_16_data_FIFO_blk[32] = 1'b0;
    assign proc_16_data_PIPO_blk[32] = 1'b0;
    assign proc_16_start_FIFO_blk[32] = 1'b0;
    assign proc_16_TLF_FIFO_blk[32] = 1'b0;
    assign proc_16_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_11_U0_ap_ready & ProcessingElement_11_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_16_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_16[32] = dl_detect_out ? proc_dep_vld_vec_16_reg[32] : (proc_16_data_FIFO_blk[32] | proc_16_data_PIPO_blk[32] | proc_16_start_FIFO_blk[32] | proc_16_TLF_FIFO_blk[32] | proc_16_input_sync_blk[32] | proc_16_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_16_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_16_reg <= proc_dep_vld_vec_16;
        end
    end
    assign in_chan_dep_vld_vec_16[0] = dep_chan_vld_0_16;
    assign in_chan_dep_data_vec_16[39 : 0] = dep_chan_data_0_16;
    assign token_in_vec_16[0] = token_0_16;
    assign in_chan_dep_vld_vec_16[1] = dep_chan_vld_1_16;
    assign in_chan_dep_data_vec_16[79 : 40] = dep_chan_data_1_16;
    assign token_in_vec_16[1] = token_1_16;
    assign in_chan_dep_vld_vec_16[2] = dep_chan_vld_3_16;
    assign in_chan_dep_data_vec_16[119 : 80] = dep_chan_data_3_16;
    assign token_in_vec_16[2] = token_3_16;
    assign in_chan_dep_vld_vec_16[3] = dep_chan_vld_6_16;
    assign in_chan_dep_data_vec_16[159 : 120] = dep_chan_data_6_16;
    assign token_in_vec_16[3] = token_6_16;
    assign in_chan_dep_vld_vec_16[4] = dep_chan_vld_7_16;
    assign in_chan_dep_data_vec_16[199 : 160] = dep_chan_data_7_16;
    assign token_in_vec_16[4] = token_7_16;
    assign in_chan_dep_vld_vec_16[5] = dep_chan_vld_8_16;
    assign in_chan_dep_data_vec_16[239 : 200] = dep_chan_data_8_16;
    assign token_in_vec_16[5] = token_8_16;
    assign in_chan_dep_vld_vec_16[6] = dep_chan_vld_9_16;
    assign in_chan_dep_data_vec_16[279 : 240] = dep_chan_data_9_16;
    assign token_in_vec_16[6] = token_9_16;
    assign in_chan_dep_vld_vec_16[7] = dep_chan_vld_10_16;
    assign in_chan_dep_data_vec_16[319 : 280] = dep_chan_data_10_16;
    assign token_in_vec_16[7] = token_10_16;
    assign in_chan_dep_vld_vec_16[8] = dep_chan_vld_11_16;
    assign in_chan_dep_data_vec_16[359 : 320] = dep_chan_data_11_16;
    assign token_in_vec_16[8] = token_11_16;
    assign in_chan_dep_vld_vec_16[9] = dep_chan_vld_12_16;
    assign in_chan_dep_data_vec_16[399 : 360] = dep_chan_data_12_16;
    assign token_in_vec_16[9] = token_12_16;
    assign in_chan_dep_vld_vec_16[10] = dep_chan_vld_13_16;
    assign in_chan_dep_data_vec_16[439 : 400] = dep_chan_data_13_16;
    assign token_in_vec_16[10] = token_13_16;
    assign in_chan_dep_vld_vec_16[11] = dep_chan_vld_14_16;
    assign in_chan_dep_data_vec_16[479 : 440] = dep_chan_data_14_16;
    assign token_in_vec_16[11] = token_14_16;
    assign in_chan_dep_vld_vec_16[12] = dep_chan_vld_15_16;
    assign in_chan_dep_data_vec_16[519 : 480] = dep_chan_data_15_16;
    assign token_in_vec_16[12] = token_15_16;
    assign in_chan_dep_vld_vec_16[13] = dep_chan_vld_17_16;
    assign in_chan_dep_data_vec_16[559 : 520] = dep_chan_data_17_16;
    assign token_in_vec_16[13] = token_17_16;
    assign in_chan_dep_vld_vec_16[14] = dep_chan_vld_18_16;
    assign in_chan_dep_data_vec_16[599 : 560] = dep_chan_data_18_16;
    assign token_in_vec_16[14] = token_18_16;
    assign in_chan_dep_vld_vec_16[15] = dep_chan_vld_19_16;
    assign in_chan_dep_data_vec_16[639 : 600] = dep_chan_data_19_16;
    assign token_in_vec_16[15] = token_19_16;
    assign in_chan_dep_vld_vec_16[16] = dep_chan_vld_20_16;
    assign in_chan_dep_data_vec_16[679 : 640] = dep_chan_data_20_16;
    assign token_in_vec_16[16] = token_20_16;
    assign in_chan_dep_vld_vec_16[17] = dep_chan_vld_21_16;
    assign in_chan_dep_data_vec_16[719 : 680] = dep_chan_data_21_16;
    assign token_in_vec_16[17] = token_21_16;
    assign in_chan_dep_vld_vec_16[18] = dep_chan_vld_22_16;
    assign in_chan_dep_data_vec_16[759 : 720] = dep_chan_data_22_16;
    assign token_in_vec_16[18] = token_22_16;
    assign in_chan_dep_vld_vec_16[19] = dep_chan_vld_23_16;
    assign in_chan_dep_data_vec_16[799 : 760] = dep_chan_data_23_16;
    assign token_in_vec_16[19] = token_23_16;
    assign in_chan_dep_vld_vec_16[20] = dep_chan_vld_24_16;
    assign in_chan_dep_data_vec_16[839 : 800] = dep_chan_data_24_16;
    assign token_in_vec_16[20] = token_24_16;
    assign in_chan_dep_vld_vec_16[21] = dep_chan_vld_25_16;
    assign in_chan_dep_data_vec_16[879 : 840] = dep_chan_data_25_16;
    assign token_in_vec_16[21] = token_25_16;
    assign in_chan_dep_vld_vec_16[22] = dep_chan_vld_26_16;
    assign in_chan_dep_data_vec_16[919 : 880] = dep_chan_data_26_16;
    assign token_in_vec_16[22] = token_26_16;
    assign in_chan_dep_vld_vec_16[23] = dep_chan_vld_27_16;
    assign in_chan_dep_data_vec_16[959 : 920] = dep_chan_data_27_16;
    assign token_in_vec_16[23] = token_27_16;
    assign in_chan_dep_vld_vec_16[24] = dep_chan_vld_28_16;
    assign in_chan_dep_data_vec_16[999 : 960] = dep_chan_data_28_16;
    assign token_in_vec_16[24] = token_28_16;
    assign in_chan_dep_vld_vec_16[25] = dep_chan_vld_29_16;
    assign in_chan_dep_data_vec_16[1039 : 1000] = dep_chan_data_29_16;
    assign token_in_vec_16[25] = token_29_16;
    assign in_chan_dep_vld_vec_16[26] = dep_chan_vld_30_16;
    assign in_chan_dep_data_vec_16[1079 : 1040] = dep_chan_data_30_16;
    assign token_in_vec_16[26] = token_30_16;
    assign in_chan_dep_vld_vec_16[27] = dep_chan_vld_31_16;
    assign in_chan_dep_data_vec_16[1119 : 1080] = dep_chan_data_31_16;
    assign token_in_vec_16[27] = token_31_16;
    assign in_chan_dep_vld_vec_16[28] = dep_chan_vld_32_16;
    assign in_chan_dep_data_vec_16[1159 : 1120] = dep_chan_data_32_16;
    assign token_in_vec_16[28] = token_32_16;
    assign in_chan_dep_vld_vec_16[29] = dep_chan_vld_33_16;
    assign in_chan_dep_data_vec_16[1199 : 1160] = dep_chan_data_33_16;
    assign token_in_vec_16[29] = token_33_16;
    assign in_chan_dep_vld_vec_16[30] = dep_chan_vld_34_16;
    assign in_chan_dep_data_vec_16[1239 : 1200] = dep_chan_data_34_16;
    assign token_in_vec_16[30] = token_34_16;
    assign in_chan_dep_vld_vec_16[31] = dep_chan_vld_35_16;
    assign in_chan_dep_data_vec_16[1279 : 1240] = dep_chan_data_35_16;
    assign token_in_vec_16[31] = token_35_16;
    assign in_chan_dep_vld_vec_16[32] = dep_chan_vld_36_16;
    assign in_chan_dep_data_vec_16[1319 : 1280] = dep_chan_data_36_16;
    assign token_in_vec_16[32] = token_36_16;
    assign dep_chan_vld_16_15 = out_chan_dep_vld_vec_16[0];
    assign dep_chan_data_16_15 = out_chan_dep_data_16;
    assign token_16_15 = token_out_vec_16[0];
    assign dep_chan_vld_16_17 = out_chan_dep_vld_vec_16[1];
    assign dep_chan_data_16_17 = out_chan_dep_data_16;
    assign token_16_17 = token_out_vec_16[1];
    assign dep_chan_vld_16_0 = out_chan_dep_vld_vec_16[2];
    assign dep_chan_data_16_0 = out_chan_dep_data_16;
    assign token_16_0 = token_out_vec_16[2];
    assign dep_chan_vld_16_1 = out_chan_dep_vld_vec_16[3];
    assign dep_chan_data_16_1 = out_chan_dep_data_16;
    assign token_16_1 = token_out_vec_16[3];
    assign dep_chan_vld_16_3 = out_chan_dep_vld_vec_16[4];
    assign dep_chan_data_16_3 = out_chan_dep_data_16;
    assign token_16_3 = token_out_vec_16[4];
    assign dep_chan_vld_16_6 = out_chan_dep_vld_vec_16[5];
    assign dep_chan_data_16_6 = out_chan_dep_data_16;
    assign token_16_6 = token_out_vec_16[5];
    assign dep_chan_vld_16_7 = out_chan_dep_vld_vec_16[6];
    assign dep_chan_data_16_7 = out_chan_dep_data_16;
    assign token_16_7 = token_out_vec_16[6];
    assign dep_chan_vld_16_8 = out_chan_dep_vld_vec_16[7];
    assign dep_chan_data_16_8 = out_chan_dep_data_16;
    assign token_16_8 = token_out_vec_16[7];
    assign dep_chan_vld_16_9 = out_chan_dep_vld_vec_16[8];
    assign dep_chan_data_16_9 = out_chan_dep_data_16;
    assign token_16_9 = token_out_vec_16[8];
    assign dep_chan_vld_16_10 = out_chan_dep_vld_vec_16[9];
    assign dep_chan_data_16_10 = out_chan_dep_data_16;
    assign token_16_10 = token_out_vec_16[9];
    assign dep_chan_vld_16_11 = out_chan_dep_vld_vec_16[10];
    assign dep_chan_data_16_11 = out_chan_dep_data_16;
    assign token_16_11 = token_out_vec_16[10];
    assign dep_chan_vld_16_12 = out_chan_dep_vld_vec_16[11];
    assign dep_chan_data_16_12 = out_chan_dep_data_16;
    assign token_16_12 = token_out_vec_16[11];
    assign dep_chan_vld_16_13 = out_chan_dep_vld_vec_16[12];
    assign dep_chan_data_16_13 = out_chan_dep_data_16;
    assign token_16_13 = token_out_vec_16[12];
    assign dep_chan_vld_16_14 = out_chan_dep_vld_vec_16[13];
    assign dep_chan_data_16_14 = out_chan_dep_data_16;
    assign token_16_14 = token_out_vec_16[13];
    assign dep_chan_vld_16_18 = out_chan_dep_vld_vec_16[14];
    assign dep_chan_data_16_18 = out_chan_dep_data_16;
    assign token_16_18 = token_out_vec_16[14];
    assign dep_chan_vld_16_19 = out_chan_dep_vld_vec_16[15];
    assign dep_chan_data_16_19 = out_chan_dep_data_16;
    assign token_16_19 = token_out_vec_16[15];
    assign dep_chan_vld_16_20 = out_chan_dep_vld_vec_16[16];
    assign dep_chan_data_16_20 = out_chan_dep_data_16;
    assign token_16_20 = token_out_vec_16[16];
    assign dep_chan_vld_16_21 = out_chan_dep_vld_vec_16[17];
    assign dep_chan_data_16_21 = out_chan_dep_data_16;
    assign token_16_21 = token_out_vec_16[17];
    assign dep_chan_vld_16_22 = out_chan_dep_vld_vec_16[18];
    assign dep_chan_data_16_22 = out_chan_dep_data_16;
    assign token_16_22 = token_out_vec_16[18];
    assign dep_chan_vld_16_23 = out_chan_dep_vld_vec_16[19];
    assign dep_chan_data_16_23 = out_chan_dep_data_16;
    assign token_16_23 = token_out_vec_16[19];
    assign dep_chan_vld_16_24 = out_chan_dep_vld_vec_16[20];
    assign dep_chan_data_16_24 = out_chan_dep_data_16;
    assign token_16_24 = token_out_vec_16[20];
    assign dep_chan_vld_16_25 = out_chan_dep_vld_vec_16[21];
    assign dep_chan_data_16_25 = out_chan_dep_data_16;
    assign token_16_25 = token_out_vec_16[21];
    assign dep_chan_vld_16_26 = out_chan_dep_vld_vec_16[22];
    assign dep_chan_data_16_26 = out_chan_dep_data_16;
    assign token_16_26 = token_out_vec_16[22];
    assign dep_chan_vld_16_27 = out_chan_dep_vld_vec_16[23];
    assign dep_chan_data_16_27 = out_chan_dep_data_16;
    assign token_16_27 = token_out_vec_16[23];
    assign dep_chan_vld_16_28 = out_chan_dep_vld_vec_16[24];
    assign dep_chan_data_16_28 = out_chan_dep_data_16;
    assign token_16_28 = token_out_vec_16[24];
    assign dep_chan_vld_16_29 = out_chan_dep_vld_vec_16[25];
    assign dep_chan_data_16_29 = out_chan_dep_data_16;
    assign token_16_29 = token_out_vec_16[25];
    assign dep_chan_vld_16_30 = out_chan_dep_vld_vec_16[26];
    assign dep_chan_data_16_30 = out_chan_dep_data_16;
    assign token_16_30 = token_out_vec_16[26];
    assign dep_chan_vld_16_31 = out_chan_dep_vld_vec_16[27];
    assign dep_chan_data_16_31 = out_chan_dep_data_16;
    assign token_16_31 = token_out_vec_16[27];
    assign dep_chan_vld_16_32 = out_chan_dep_vld_vec_16[28];
    assign dep_chan_data_16_32 = out_chan_dep_data_16;
    assign token_16_32 = token_out_vec_16[28];
    assign dep_chan_vld_16_33 = out_chan_dep_vld_vec_16[29];
    assign dep_chan_data_16_33 = out_chan_dep_data_16;
    assign token_16_33 = token_out_vec_16[29];
    assign dep_chan_vld_16_34 = out_chan_dep_vld_vec_16[30];
    assign dep_chan_data_16_34 = out_chan_dep_data_16;
    assign token_16_34 = token_out_vec_16[30];
    assign dep_chan_vld_16_35 = out_chan_dep_vld_vec_16[31];
    assign dep_chan_data_16_35 = out_chan_dep_data_16;
    assign token_16_35 = token_out_vec_16[31];
    assign dep_chan_vld_16_36 = out_chan_dep_vld_vec_16[32];
    assign dep_chan_data_16_36 = out_chan_dep_data_16;
    assign token_16_36 = token_out_vec_16[32];

    // Process: ProcessingElement_12_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 17, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_17 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_17),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_17),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_17),
        .token_in_vec(token_in_vec_17),
        .dl_detect_in(dl_detect_out),
        .origin(origin[17]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_17),
        .out_chan_dep_data(out_chan_dep_data_17),
        .token_out_vec(token_out_vec_17),
        .dl_detect_out(dl_in_vec[17]));

    assign proc_17_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_11_blk_n) | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_11_blk_n) | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_WriteC_Flattened_fu_179.cPipes_11_blk_n);
    assign proc_17_data_PIPO_blk[0] = 1'b0;
    assign proc_17_start_FIFO_blk[0] = 1'b0;
    assign proc_17_TLF_FIFO_blk[0] = 1'b0;
    assign proc_17_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_17_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_17[0] = dl_detect_out ? proc_dep_vld_vec_17_reg[0] : (proc_17_data_FIFO_blk[0] | proc_17_data_PIPO_blk[0] | proc_17_start_FIFO_blk[0] | proc_17_TLF_FIFO_blk[0] | proc_17_input_sync_blk[0] | proc_17_output_sync_blk[0]);
    assign proc_17_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_12_blk_n) | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_12_blk_n) | (~ProcessingElement_12_U0.grp_ProcessingElement_12_Pipeline_WriteC_Flattened_fu_179.cPipes_12_blk_n);
    assign proc_17_data_PIPO_blk[1] = 1'b0;
    assign proc_17_start_FIFO_blk[1] = 1'b0;
    assign proc_17_TLF_FIFO_blk[1] = 1'b0;
    assign proc_17_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_17_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_17[1] = dl_detect_out ? proc_dep_vld_vec_17_reg[1] : (proc_17_data_FIFO_blk[1] | proc_17_data_PIPO_blk[1] | proc_17_start_FIFO_blk[1] | proc_17_TLF_FIFO_blk[1] | proc_17_input_sync_blk[1] | proc_17_output_sync_blk[1]);
    assign proc_17_data_FIFO_blk[2] = 1'b0;
    assign proc_17_data_PIPO_blk[2] = 1'b0;
    assign proc_17_start_FIFO_blk[2] = 1'b0;
    assign proc_17_TLF_FIFO_blk[2] = 1'b0;
    assign proc_17_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_17_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_17[2] = dl_detect_out ? proc_dep_vld_vec_17_reg[2] : (proc_17_data_FIFO_blk[2] | proc_17_data_PIPO_blk[2] | proc_17_start_FIFO_blk[2] | proc_17_TLF_FIFO_blk[2] | proc_17_input_sync_blk[2] | proc_17_output_sync_blk[2]);
    assign proc_17_data_FIFO_blk[3] = 1'b0;
    assign proc_17_data_PIPO_blk[3] = 1'b0;
    assign proc_17_start_FIFO_blk[3] = 1'b0;
    assign proc_17_TLF_FIFO_blk[3] = 1'b0;
    assign proc_17_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_17_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_17[3] = dl_detect_out ? proc_dep_vld_vec_17_reg[3] : (proc_17_data_FIFO_blk[3] | proc_17_data_PIPO_blk[3] | proc_17_start_FIFO_blk[3] | proc_17_TLF_FIFO_blk[3] | proc_17_input_sync_blk[3] | proc_17_output_sync_blk[3]);
    assign proc_17_data_FIFO_blk[4] = 1'b0;
    assign proc_17_data_PIPO_blk[4] = 1'b0;
    assign proc_17_start_FIFO_blk[4] = 1'b0;
    assign proc_17_TLF_FIFO_blk[4] = 1'b0;
    assign proc_17_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_17_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_17[4] = dl_detect_out ? proc_dep_vld_vec_17_reg[4] : (proc_17_data_FIFO_blk[4] | proc_17_data_PIPO_blk[4] | proc_17_start_FIFO_blk[4] | proc_17_TLF_FIFO_blk[4] | proc_17_input_sync_blk[4] | proc_17_output_sync_blk[4]);
    assign proc_17_data_FIFO_blk[5] = 1'b0;
    assign proc_17_data_PIPO_blk[5] = 1'b0;
    assign proc_17_start_FIFO_blk[5] = 1'b0;
    assign proc_17_TLF_FIFO_blk[5] = 1'b0;
    assign proc_17_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_17_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_17[5] = dl_detect_out ? proc_dep_vld_vec_17_reg[5] : (proc_17_data_FIFO_blk[5] | proc_17_data_PIPO_blk[5] | proc_17_start_FIFO_blk[5] | proc_17_TLF_FIFO_blk[5] | proc_17_input_sync_blk[5] | proc_17_output_sync_blk[5]);
    assign proc_17_data_FIFO_blk[6] = 1'b0;
    assign proc_17_data_PIPO_blk[6] = 1'b0;
    assign proc_17_start_FIFO_blk[6] = 1'b0;
    assign proc_17_TLF_FIFO_blk[6] = 1'b0;
    assign proc_17_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_17_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_17[6] = dl_detect_out ? proc_dep_vld_vec_17_reg[6] : (proc_17_data_FIFO_blk[6] | proc_17_data_PIPO_blk[6] | proc_17_start_FIFO_blk[6] | proc_17_TLF_FIFO_blk[6] | proc_17_input_sync_blk[6] | proc_17_output_sync_blk[6]);
    assign proc_17_data_FIFO_blk[7] = 1'b0;
    assign proc_17_data_PIPO_blk[7] = 1'b0;
    assign proc_17_start_FIFO_blk[7] = 1'b0;
    assign proc_17_TLF_FIFO_blk[7] = 1'b0;
    assign proc_17_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_17_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_17[7] = dl_detect_out ? proc_dep_vld_vec_17_reg[7] : (proc_17_data_FIFO_blk[7] | proc_17_data_PIPO_blk[7] | proc_17_start_FIFO_blk[7] | proc_17_TLF_FIFO_blk[7] | proc_17_input_sync_blk[7] | proc_17_output_sync_blk[7]);
    assign proc_17_data_FIFO_blk[8] = 1'b0;
    assign proc_17_data_PIPO_blk[8] = 1'b0;
    assign proc_17_start_FIFO_blk[8] = 1'b0;
    assign proc_17_TLF_FIFO_blk[8] = 1'b0;
    assign proc_17_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_17_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_17[8] = dl_detect_out ? proc_dep_vld_vec_17_reg[8] : (proc_17_data_FIFO_blk[8] | proc_17_data_PIPO_blk[8] | proc_17_start_FIFO_blk[8] | proc_17_TLF_FIFO_blk[8] | proc_17_input_sync_blk[8] | proc_17_output_sync_blk[8]);
    assign proc_17_data_FIFO_blk[9] = 1'b0;
    assign proc_17_data_PIPO_blk[9] = 1'b0;
    assign proc_17_start_FIFO_blk[9] = 1'b0;
    assign proc_17_TLF_FIFO_blk[9] = 1'b0;
    assign proc_17_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_17_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_17[9] = dl_detect_out ? proc_dep_vld_vec_17_reg[9] : (proc_17_data_FIFO_blk[9] | proc_17_data_PIPO_blk[9] | proc_17_start_FIFO_blk[9] | proc_17_TLF_FIFO_blk[9] | proc_17_input_sync_blk[9] | proc_17_output_sync_blk[9]);
    assign proc_17_data_FIFO_blk[10] = 1'b0;
    assign proc_17_data_PIPO_blk[10] = 1'b0;
    assign proc_17_start_FIFO_blk[10] = 1'b0;
    assign proc_17_TLF_FIFO_blk[10] = 1'b0;
    assign proc_17_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_17_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_17[10] = dl_detect_out ? proc_dep_vld_vec_17_reg[10] : (proc_17_data_FIFO_blk[10] | proc_17_data_PIPO_blk[10] | proc_17_start_FIFO_blk[10] | proc_17_TLF_FIFO_blk[10] | proc_17_input_sync_blk[10] | proc_17_output_sync_blk[10]);
    assign proc_17_data_FIFO_blk[11] = 1'b0;
    assign proc_17_data_PIPO_blk[11] = 1'b0;
    assign proc_17_start_FIFO_blk[11] = 1'b0;
    assign proc_17_TLF_FIFO_blk[11] = 1'b0;
    assign proc_17_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_17_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_17[11] = dl_detect_out ? proc_dep_vld_vec_17_reg[11] : (proc_17_data_FIFO_blk[11] | proc_17_data_PIPO_blk[11] | proc_17_start_FIFO_blk[11] | proc_17_TLF_FIFO_blk[11] | proc_17_input_sync_blk[11] | proc_17_output_sync_blk[11]);
    assign proc_17_data_FIFO_blk[12] = 1'b0;
    assign proc_17_data_PIPO_blk[12] = 1'b0;
    assign proc_17_start_FIFO_blk[12] = 1'b0;
    assign proc_17_TLF_FIFO_blk[12] = 1'b0;
    assign proc_17_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_17_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_17[12] = dl_detect_out ? proc_dep_vld_vec_17_reg[12] : (proc_17_data_FIFO_blk[12] | proc_17_data_PIPO_blk[12] | proc_17_start_FIFO_blk[12] | proc_17_TLF_FIFO_blk[12] | proc_17_input_sync_blk[12] | proc_17_output_sync_blk[12]);
    assign proc_17_data_FIFO_blk[13] = 1'b0;
    assign proc_17_data_PIPO_blk[13] = 1'b0;
    assign proc_17_start_FIFO_blk[13] = 1'b0;
    assign proc_17_TLF_FIFO_blk[13] = 1'b0;
    assign proc_17_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_17_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_17[13] = dl_detect_out ? proc_dep_vld_vec_17_reg[13] : (proc_17_data_FIFO_blk[13] | proc_17_data_PIPO_blk[13] | proc_17_start_FIFO_blk[13] | proc_17_TLF_FIFO_blk[13] | proc_17_input_sync_blk[13] | proc_17_output_sync_blk[13]);
    assign proc_17_data_FIFO_blk[14] = 1'b0;
    assign proc_17_data_PIPO_blk[14] = 1'b0;
    assign proc_17_start_FIFO_blk[14] = 1'b0;
    assign proc_17_TLF_FIFO_blk[14] = 1'b0;
    assign proc_17_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_17_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_17[14] = dl_detect_out ? proc_dep_vld_vec_17_reg[14] : (proc_17_data_FIFO_blk[14] | proc_17_data_PIPO_blk[14] | proc_17_start_FIFO_blk[14] | proc_17_TLF_FIFO_blk[14] | proc_17_input_sync_blk[14] | proc_17_output_sync_blk[14]);
    assign proc_17_data_FIFO_blk[15] = 1'b0;
    assign proc_17_data_PIPO_blk[15] = 1'b0;
    assign proc_17_start_FIFO_blk[15] = 1'b0;
    assign proc_17_TLF_FIFO_blk[15] = 1'b0;
    assign proc_17_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_17_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_17[15] = dl_detect_out ? proc_dep_vld_vec_17_reg[15] : (proc_17_data_FIFO_blk[15] | proc_17_data_PIPO_blk[15] | proc_17_start_FIFO_blk[15] | proc_17_TLF_FIFO_blk[15] | proc_17_input_sync_blk[15] | proc_17_output_sync_blk[15]);
    assign proc_17_data_FIFO_blk[16] = 1'b0;
    assign proc_17_data_PIPO_blk[16] = 1'b0;
    assign proc_17_start_FIFO_blk[16] = 1'b0;
    assign proc_17_TLF_FIFO_blk[16] = 1'b0;
    assign proc_17_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_17_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_17[16] = dl_detect_out ? proc_dep_vld_vec_17_reg[16] : (proc_17_data_FIFO_blk[16] | proc_17_data_PIPO_blk[16] | proc_17_start_FIFO_blk[16] | proc_17_TLF_FIFO_blk[16] | proc_17_input_sync_blk[16] | proc_17_output_sync_blk[16]);
    assign proc_17_data_FIFO_blk[17] = 1'b0;
    assign proc_17_data_PIPO_blk[17] = 1'b0;
    assign proc_17_start_FIFO_blk[17] = 1'b0;
    assign proc_17_TLF_FIFO_blk[17] = 1'b0;
    assign proc_17_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_17_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_17[17] = dl_detect_out ? proc_dep_vld_vec_17_reg[17] : (proc_17_data_FIFO_blk[17] | proc_17_data_PIPO_blk[17] | proc_17_start_FIFO_blk[17] | proc_17_TLF_FIFO_blk[17] | proc_17_input_sync_blk[17] | proc_17_output_sync_blk[17]);
    assign proc_17_data_FIFO_blk[18] = 1'b0;
    assign proc_17_data_PIPO_blk[18] = 1'b0;
    assign proc_17_start_FIFO_blk[18] = 1'b0;
    assign proc_17_TLF_FIFO_blk[18] = 1'b0;
    assign proc_17_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_17_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_17[18] = dl_detect_out ? proc_dep_vld_vec_17_reg[18] : (proc_17_data_FIFO_blk[18] | proc_17_data_PIPO_blk[18] | proc_17_start_FIFO_blk[18] | proc_17_TLF_FIFO_blk[18] | proc_17_input_sync_blk[18] | proc_17_output_sync_blk[18]);
    assign proc_17_data_FIFO_blk[19] = 1'b0;
    assign proc_17_data_PIPO_blk[19] = 1'b0;
    assign proc_17_start_FIFO_blk[19] = 1'b0;
    assign proc_17_TLF_FIFO_blk[19] = 1'b0;
    assign proc_17_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_17_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_17[19] = dl_detect_out ? proc_dep_vld_vec_17_reg[19] : (proc_17_data_FIFO_blk[19] | proc_17_data_PIPO_blk[19] | proc_17_start_FIFO_blk[19] | proc_17_TLF_FIFO_blk[19] | proc_17_input_sync_blk[19] | proc_17_output_sync_blk[19]);
    assign proc_17_data_FIFO_blk[20] = 1'b0;
    assign proc_17_data_PIPO_blk[20] = 1'b0;
    assign proc_17_start_FIFO_blk[20] = 1'b0;
    assign proc_17_TLF_FIFO_blk[20] = 1'b0;
    assign proc_17_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_17_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_17[20] = dl_detect_out ? proc_dep_vld_vec_17_reg[20] : (proc_17_data_FIFO_blk[20] | proc_17_data_PIPO_blk[20] | proc_17_start_FIFO_blk[20] | proc_17_TLF_FIFO_blk[20] | proc_17_input_sync_blk[20] | proc_17_output_sync_blk[20]);
    assign proc_17_data_FIFO_blk[21] = 1'b0;
    assign proc_17_data_PIPO_blk[21] = 1'b0;
    assign proc_17_start_FIFO_blk[21] = 1'b0;
    assign proc_17_TLF_FIFO_blk[21] = 1'b0;
    assign proc_17_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_17_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_17[21] = dl_detect_out ? proc_dep_vld_vec_17_reg[21] : (proc_17_data_FIFO_blk[21] | proc_17_data_PIPO_blk[21] | proc_17_start_FIFO_blk[21] | proc_17_TLF_FIFO_blk[21] | proc_17_input_sync_blk[21] | proc_17_output_sync_blk[21]);
    assign proc_17_data_FIFO_blk[22] = 1'b0;
    assign proc_17_data_PIPO_blk[22] = 1'b0;
    assign proc_17_start_FIFO_blk[22] = 1'b0;
    assign proc_17_TLF_FIFO_blk[22] = 1'b0;
    assign proc_17_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_17_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_17[22] = dl_detect_out ? proc_dep_vld_vec_17_reg[22] : (proc_17_data_FIFO_blk[22] | proc_17_data_PIPO_blk[22] | proc_17_start_FIFO_blk[22] | proc_17_TLF_FIFO_blk[22] | proc_17_input_sync_blk[22] | proc_17_output_sync_blk[22]);
    assign proc_17_data_FIFO_blk[23] = 1'b0;
    assign proc_17_data_PIPO_blk[23] = 1'b0;
    assign proc_17_start_FIFO_blk[23] = 1'b0;
    assign proc_17_TLF_FIFO_blk[23] = 1'b0;
    assign proc_17_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_17_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_17[23] = dl_detect_out ? proc_dep_vld_vec_17_reg[23] : (proc_17_data_FIFO_blk[23] | proc_17_data_PIPO_blk[23] | proc_17_start_FIFO_blk[23] | proc_17_TLF_FIFO_blk[23] | proc_17_input_sync_blk[23] | proc_17_output_sync_blk[23]);
    assign proc_17_data_FIFO_blk[24] = 1'b0;
    assign proc_17_data_PIPO_blk[24] = 1'b0;
    assign proc_17_start_FIFO_blk[24] = 1'b0;
    assign proc_17_TLF_FIFO_blk[24] = 1'b0;
    assign proc_17_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_17_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_17[24] = dl_detect_out ? proc_dep_vld_vec_17_reg[24] : (proc_17_data_FIFO_blk[24] | proc_17_data_PIPO_blk[24] | proc_17_start_FIFO_blk[24] | proc_17_TLF_FIFO_blk[24] | proc_17_input_sync_blk[24] | proc_17_output_sync_blk[24]);
    assign proc_17_data_FIFO_blk[25] = 1'b0;
    assign proc_17_data_PIPO_blk[25] = 1'b0;
    assign proc_17_start_FIFO_blk[25] = 1'b0;
    assign proc_17_TLF_FIFO_blk[25] = 1'b0;
    assign proc_17_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_17_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_17[25] = dl_detect_out ? proc_dep_vld_vec_17_reg[25] : (proc_17_data_FIFO_blk[25] | proc_17_data_PIPO_blk[25] | proc_17_start_FIFO_blk[25] | proc_17_TLF_FIFO_blk[25] | proc_17_input_sync_blk[25] | proc_17_output_sync_blk[25]);
    assign proc_17_data_FIFO_blk[26] = 1'b0;
    assign proc_17_data_PIPO_blk[26] = 1'b0;
    assign proc_17_start_FIFO_blk[26] = 1'b0;
    assign proc_17_TLF_FIFO_blk[26] = 1'b0;
    assign proc_17_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_17_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_17[26] = dl_detect_out ? proc_dep_vld_vec_17_reg[26] : (proc_17_data_FIFO_blk[26] | proc_17_data_PIPO_blk[26] | proc_17_start_FIFO_blk[26] | proc_17_TLF_FIFO_blk[26] | proc_17_input_sync_blk[26] | proc_17_output_sync_blk[26]);
    assign proc_17_data_FIFO_blk[27] = 1'b0;
    assign proc_17_data_PIPO_blk[27] = 1'b0;
    assign proc_17_start_FIFO_blk[27] = 1'b0;
    assign proc_17_TLF_FIFO_blk[27] = 1'b0;
    assign proc_17_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_17_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_17[27] = dl_detect_out ? proc_dep_vld_vec_17_reg[27] : (proc_17_data_FIFO_blk[27] | proc_17_data_PIPO_blk[27] | proc_17_start_FIFO_blk[27] | proc_17_TLF_FIFO_blk[27] | proc_17_input_sync_blk[27] | proc_17_output_sync_blk[27]);
    assign proc_17_data_FIFO_blk[28] = 1'b0;
    assign proc_17_data_PIPO_blk[28] = 1'b0;
    assign proc_17_start_FIFO_blk[28] = 1'b0;
    assign proc_17_TLF_FIFO_blk[28] = 1'b0;
    assign proc_17_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_17_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_17[28] = dl_detect_out ? proc_dep_vld_vec_17_reg[28] : (proc_17_data_FIFO_blk[28] | proc_17_data_PIPO_blk[28] | proc_17_start_FIFO_blk[28] | proc_17_TLF_FIFO_blk[28] | proc_17_input_sync_blk[28] | proc_17_output_sync_blk[28]);
    assign proc_17_data_FIFO_blk[29] = 1'b0;
    assign proc_17_data_PIPO_blk[29] = 1'b0;
    assign proc_17_start_FIFO_blk[29] = 1'b0;
    assign proc_17_TLF_FIFO_blk[29] = 1'b0;
    assign proc_17_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_17_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_17[29] = dl_detect_out ? proc_dep_vld_vec_17_reg[29] : (proc_17_data_FIFO_blk[29] | proc_17_data_PIPO_blk[29] | proc_17_start_FIFO_blk[29] | proc_17_TLF_FIFO_blk[29] | proc_17_input_sync_blk[29] | proc_17_output_sync_blk[29]);
    assign proc_17_data_FIFO_blk[30] = 1'b0;
    assign proc_17_data_PIPO_blk[30] = 1'b0;
    assign proc_17_start_FIFO_blk[30] = 1'b0;
    assign proc_17_TLF_FIFO_blk[30] = 1'b0;
    assign proc_17_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_17_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_17[30] = dl_detect_out ? proc_dep_vld_vec_17_reg[30] : (proc_17_data_FIFO_blk[30] | proc_17_data_PIPO_blk[30] | proc_17_start_FIFO_blk[30] | proc_17_TLF_FIFO_blk[30] | proc_17_input_sync_blk[30] | proc_17_output_sync_blk[30]);
    assign proc_17_data_FIFO_blk[31] = 1'b0;
    assign proc_17_data_PIPO_blk[31] = 1'b0;
    assign proc_17_start_FIFO_blk[31] = 1'b0;
    assign proc_17_TLF_FIFO_blk[31] = 1'b0;
    assign proc_17_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_17_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_17[31] = dl_detect_out ? proc_dep_vld_vec_17_reg[31] : (proc_17_data_FIFO_blk[31] | proc_17_data_PIPO_blk[31] | proc_17_start_FIFO_blk[31] | proc_17_TLF_FIFO_blk[31] | proc_17_input_sync_blk[31] | proc_17_output_sync_blk[31]);
    assign proc_17_data_FIFO_blk[32] = 1'b0;
    assign proc_17_data_PIPO_blk[32] = 1'b0;
    assign proc_17_start_FIFO_blk[32] = 1'b0;
    assign proc_17_TLF_FIFO_blk[32] = 1'b0;
    assign proc_17_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_12_U0_ap_ready & ProcessingElement_12_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_17_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_17[32] = dl_detect_out ? proc_dep_vld_vec_17_reg[32] : (proc_17_data_FIFO_blk[32] | proc_17_data_PIPO_blk[32] | proc_17_start_FIFO_blk[32] | proc_17_TLF_FIFO_blk[32] | proc_17_input_sync_blk[32] | proc_17_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_17_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_17_reg <= proc_dep_vld_vec_17;
        end
    end
    assign in_chan_dep_vld_vec_17[0] = dep_chan_vld_0_17;
    assign in_chan_dep_data_vec_17[39 : 0] = dep_chan_data_0_17;
    assign token_in_vec_17[0] = token_0_17;
    assign in_chan_dep_vld_vec_17[1] = dep_chan_vld_1_17;
    assign in_chan_dep_data_vec_17[79 : 40] = dep_chan_data_1_17;
    assign token_in_vec_17[1] = token_1_17;
    assign in_chan_dep_vld_vec_17[2] = dep_chan_vld_3_17;
    assign in_chan_dep_data_vec_17[119 : 80] = dep_chan_data_3_17;
    assign token_in_vec_17[2] = token_3_17;
    assign in_chan_dep_vld_vec_17[3] = dep_chan_vld_6_17;
    assign in_chan_dep_data_vec_17[159 : 120] = dep_chan_data_6_17;
    assign token_in_vec_17[3] = token_6_17;
    assign in_chan_dep_vld_vec_17[4] = dep_chan_vld_7_17;
    assign in_chan_dep_data_vec_17[199 : 160] = dep_chan_data_7_17;
    assign token_in_vec_17[4] = token_7_17;
    assign in_chan_dep_vld_vec_17[5] = dep_chan_vld_8_17;
    assign in_chan_dep_data_vec_17[239 : 200] = dep_chan_data_8_17;
    assign token_in_vec_17[5] = token_8_17;
    assign in_chan_dep_vld_vec_17[6] = dep_chan_vld_9_17;
    assign in_chan_dep_data_vec_17[279 : 240] = dep_chan_data_9_17;
    assign token_in_vec_17[6] = token_9_17;
    assign in_chan_dep_vld_vec_17[7] = dep_chan_vld_10_17;
    assign in_chan_dep_data_vec_17[319 : 280] = dep_chan_data_10_17;
    assign token_in_vec_17[7] = token_10_17;
    assign in_chan_dep_vld_vec_17[8] = dep_chan_vld_11_17;
    assign in_chan_dep_data_vec_17[359 : 320] = dep_chan_data_11_17;
    assign token_in_vec_17[8] = token_11_17;
    assign in_chan_dep_vld_vec_17[9] = dep_chan_vld_12_17;
    assign in_chan_dep_data_vec_17[399 : 360] = dep_chan_data_12_17;
    assign token_in_vec_17[9] = token_12_17;
    assign in_chan_dep_vld_vec_17[10] = dep_chan_vld_13_17;
    assign in_chan_dep_data_vec_17[439 : 400] = dep_chan_data_13_17;
    assign token_in_vec_17[10] = token_13_17;
    assign in_chan_dep_vld_vec_17[11] = dep_chan_vld_14_17;
    assign in_chan_dep_data_vec_17[479 : 440] = dep_chan_data_14_17;
    assign token_in_vec_17[11] = token_14_17;
    assign in_chan_dep_vld_vec_17[12] = dep_chan_vld_15_17;
    assign in_chan_dep_data_vec_17[519 : 480] = dep_chan_data_15_17;
    assign token_in_vec_17[12] = token_15_17;
    assign in_chan_dep_vld_vec_17[13] = dep_chan_vld_16_17;
    assign in_chan_dep_data_vec_17[559 : 520] = dep_chan_data_16_17;
    assign token_in_vec_17[13] = token_16_17;
    assign in_chan_dep_vld_vec_17[14] = dep_chan_vld_18_17;
    assign in_chan_dep_data_vec_17[599 : 560] = dep_chan_data_18_17;
    assign token_in_vec_17[14] = token_18_17;
    assign in_chan_dep_vld_vec_17[15] = dep_chan_vld_19_17;
    assign in_chan_dep_data_vec_17[639 : 600] = dep_chan_data_19_17;
    assign token_in_vec_17[15] = token_19_17;
    assign in_chan_dep_vld_vec_17[16] = dep_chan_vld_20_17;
    assign in_chan_dep_data_vec_17[679 : 640] = dep_chan_data_20_17;
    assign token_in_vec_17[16] = token_20_17;
    assign in_chan_dep_vld_vec_17[17] = dep_chan_vld_21_17;
    assign in_chan_dep_data_vec_17[719 : 680] = dep_chan_data_21_17;
    assign token_in_vec_17[17] = token_21_17;
    assign in_chan_dep_vld_vec_17[18] = dep_chan_vld_22_17;
    assign in_chan_dep_data_vec_17[759 : 720] = dep_chan_data_22_17;
    assign token_in_vec_17[18] = token_22_17;
    assign in_chan_dep_vld_vec_17[19] = dep_chan_vld_23_17;
    assign in_chan_dep_data_vec_17[799 : 760] = dep_chan_data_23_17;
    assign token_in_vec_17[19] = token_23_17;
    assign in_chan_dep_vld_vec_17[20] = dep_chan_vld_24_17;
    assign in_chan_dep_data_vec_17[839 : 800] = dep_chan_data_24_17;
    assign token_in_vec_17[20] = token_24_17;
    assign in_chan_dep_vld_vec_17[21] = dep_chan_vld_25_17;
    assign in_chan_dep_data_vec_17[879 : 840] = dep_chan_data_25_17;
    assign token_in_vec_17[21] = token_25_17;
    assign in_chan_dep_vld_vec_17[22] = dep_chan_vld_26_17;
    assign in_chan_dep_data_vec_17[919 : 880] = dep_chan_data_26_17;
    assign token_in_vec_17[22] = token_26_17;
    assign in_chan_dep_vld_vec_17[23] = dep_chan_vld_27_17;
    assign in_chan_dep_data_vec_17[959 : 920] = dep_chan_data_27_17;
    assign token_in_vec_17[23] = token_27_17;
    assign in_chan_dep_vld_vec_17[24] = dep_chan_vld_28_17;
    assign in_chan_dep_data_vec_17[999 : 960] = dep_chan_data_28_17;
    assign token_in_vec_17[24] = token_28_17;
    assign in_chan_dep_vld_vec_17[25] = dep_chan_vld_29_17;
    assign in_chan_dep_data_vec_17[1039 : 1000] = dep_chan_data_29_17;
    assign token_in_vec_17[25] = token_29_17;
    assign in_chan_dep_vld_vec_17[26] = dep_chan_vld_30_17;
    assign in_chan_dep_data_vec_17[1079 : 1040] = dep_chan_data_30_17;
    assign token_in_vec_17[26] = token_30_17;
    assign in_chan_dep_vld_vec_17[27] = dep_chan_vld_31_17;
    assign in_chan_dep_data_vec_17[1119 : 1080] = dep_chan_data_31_17;
    assign token_in_vec_17[27] = token_31_17;
    assign in_chan_dep_vld_vec_17[28] = dep_chan_vld_32_17;
    assign in_chan_dep_data_vec_17[1159 : 1120] = dep_chan_data_32_17;
    assign token_in_vec_17[28] = token_32_17;
    assign in_chan_dep_vld_vec_17[29] = dep_chan_vld_33_17;
    assign in_chan_dep_data_vec_17[1199 : 1160] = dep_chan_data_33_17;
    assign token_in_vec_17[29] = token_33_17;
    assign in_chan_dep_vld_vec_17[30] = dep_chan_vld_34_17;
    assign in_chan_dep_data_vec_17[1239 : 1200] = dep_chan_data_34_17;
    assign token_in_vec_17[30] = token_34_17;
    assign in_chan_dep_vld_vec_17[31] = dep_chan_vld_35_17;
    assign in_chan_dep_data_vec_17[1279 : 1240] = dep_chan_data_35_17;
    assign token_in_vec_17[31] = token_35_17;
    assign in_chan_dep_vld_vec_17[32] = dep_chan_vld_36_17;
    assign in_chan_dep_data_vec_17[1319 : 1280] = dep_chan_data_36_17;
    assign token_in_vec_17[32] = token_36_17;
    assign dep_chan_vld_17_16 = out_chan_dep_vld_vec_17[0];
    assign dep_chan_data_17_16 = out_chan_dep_data_17;
    assign token_17_16 = token_out_vec_17[0];
    assign dep_chan_vld_17_18 = out_chan_dep_vld_vec_17[1];
    assign dep_chan_data_17_18 = out_chan_dep_data_17;
    assign token_17_18 = token_out_vec_17[1];
    assign dep_chan_vld_17_0 = out_chan_dep_vld_vec_17[2];
    assign dep_chan_data_17_0 = out_chan_dep_data_17;
    assign token_17_0 = token_out_vec_17[2];
    assign dep_chan_vld_17_1 = out_chan_dep_vld_vec_17[3];
    assign dep_chan_data_17_1 = out_chan_dep_data_17;
    assign token_17_1 = token_out_vec_17[3];
    assign dep_chan_vld_17_3 = out_chan_dep_vld_vec_17[4];
    assign dep_chan_data_17_3 = out_chan_dep_data_17;
    assign token_17_3 = token_out_vec_17[4];
    assign dep_chan_vld_17_6 = out_chan_dep_vld_vec_17[5];
    assign dep_chan_data_17_6 = out_chan_dep_data_17;
    assign token_17_6 = token_out_vec_17[5];
    assign dep_chan_vld_17_7 = out_chan_dep_vld_vec_17[6];
    assign dep_chan_data_17_7 = out_chan_dep_data_17;
    assign token_17_7 = token_out_vec_17[6];
    assign dep_chan_vld_17_8 = out_chan_dep_vld_vec_17[7];
    assign dep_chan_data_17_8 = out_chan_dep_data_17;
    assign token_17_8 = token_out_vec_17[7];
    assign dep_chan_vld_17_9 = out_chan_dep_vld_vec_17[8];
    assign dep_chan_data_17_9 = out_chan_dep_data_17;
    assign token_17_9 = token_out_vec_17[8];
    assign dep_chan_vld_17_10 = out_chan_dep_vld_vec_17[9];
    assign dep_chan_data_17_10 = out_chan_dep_data_17;
    assign token_17_10 = token_out_vec_17[9];
    assign dep_chan_vld_17_11 = out_chan_dep_vld_vec_17[10];
    assign dep_chan_data_17_11 = out_chan_dep_data_17;
    assign token_17_11 = token_out_vec_17[10];
    assign dep_chan_vld_17_12 = out_chan_dep_vld_vec_17[11];
    assign dep_chan_data_17_12 = out_chan_dep_data_17;
    assign token_17_12 = token_out_vec_17[11];
    assign dep_chan_vld_17_13 = out_chan_dep_vld_vec_17[12];
    assign dep_chan_data_17_13 = out_chan_dep_data_17;
    assign token_17_13 = token_out_vec_17[12];
    assign dep_chan_vld_17_14 = out_chan_dep_vld_vec_17[13];
    assign dep_chan_data_17_14 = out_chan_dep_data_17;
    assign token_17_14 = token_out_vec_17[13];
    assign dep_chan_vld_17_15 = out_chan_dep_vld_vec_17[14];
    assign dep_chan_data_17_15 = out_chan_dep_data_17;
    assign token_17_15 = token_out_vec_17[14];
    assign dep_chan_vld_17_19 = out_chan_dep_vld_vec_17[15];
    assign dep_chan_data_17_19 = out_chan_dep_data_17;
    assign token_17_19 = token_out_vec_17[15];
    assign dep_chan_vld_17_20 = out_chan_dep_vld_vec_17[16];
    assign dep_chan_data_17_20 = out_chan_dep_data_17;
    assign token_17_20 = token_out_vec_17[16];
    assign dep_chan_vld_17_21 = out_chan_dep_vld_vec_17[17];
    assign dep_chan_data_17_21 = out_chan_dep_data_17;
    assign token_17_21 = token_out_vec_17[17];
    assign dep_chan_vld_17_22 = out_chan_dep_vld_vec_17[18];
    assign dep_chan_data_17_22 = out_chan_dep_data_17;
    assign token_17_22 = token_out_vec_17[18];
    assign dep_chan_vld_17_23 = out_chan_dep_vld_vec_17[19];
    assign dep_chan_data_17_23 = out_chan_dep_data_17;
    assign token_17_23 = token_out_vec_17[19];
    assign dep_chan_vld_17_24 = out_chan_dep_vld_vec_17[20];
    assign dep_chan_data_17_24 = out_chan_dep_data_17;
    assign token_17_24 = token_out_vec_17[20];
    assign dep_chan_vld_17_25 = out_chan_dep_vld_vec_17[21];
    assign dep_chan_data_17_25 = out_chan_dep_data_17;
    assign token_17_25 = token_out_vec_17[21];
    assign dep_chan_vld_17_26 = out_chan_dep_vld_vec_17[22];
    assign dep_chan_data_17_26 = out_chan_dep_data_17;
    assign token_17_26 = token_out_vec_17[22];
    assign dep_chan_vld_17_27 = out_chan_dep_vld_vec_17[23];
    assign dep_chan_data_17_27 = out_chan_dep_data_17;
    assign token_17_27 = token_out_vec_17[23];
    assign dep_chan_vld_17_28 = out_chan_dep_vld_vec_17[24];
    assign dep_chan_data_17_28 = out_chan_dep_data_17;
    assign token_17_28 = token_out_vec_17[24];
    assign dep_chan_vld_17_29 = out_chan_dep_vld_vec_17[25];
    assign dep_chan_data_17_29 = out_chan_dep_data_17;
    assign token_17_29 = token_out_vec_17[25];
    assign dep_chan_vld_17_30 = out_chan_dep_vld_vec_17[26];
    assign dep_chan_data_17_30 = out_chan_dep_data_17;
    assign token_17_30 = token_out_vec_17[26];
    assign dep_chan_vld_17_31 = out_chan_dep_vld_vec_17[27];
    assign dep_chan_data_17_31 = out_chan_dep_data_17;
    assign token_17_31 = token_out_vec_17[27];
    assign dep_chan_vld_17_32 = out_chan_dep_vld_vec_17[28];
    assign dep_chan_data_17_32 = out_chan_dep_data_17;
    assign token_17_32 = token_out_vec_17[28];
    assign dep_chan_vld_17_33 = out_chan_dep_vld_vec_17[29];
    assign dep_chan_data_17_33 = out_chan_dep_data_17;
    assign token_17_33 = token_out_vec_17[29];
    assign dep_chan_vld_17_34 = out_chan_dep_vld_vec_17[30];
    assign dep_chan_data_17_34 = out_chan_dep_data_17;
    assign token_17_34 = token_out_vec_17[30];
    assign dep_chan_vld_17_35 = out_chan_dep_vld_vec_17[31];
    assign dep_chan_data_17_35 = out_chan_dep_data_17;
    assign token_17_35 = token_out_vec_17[31];
    assign dep_chan_vld_17_36 = out_chan_dep_vld_vec_17[32];
    assign dep_chan_data_17_36 = out_chan_dep_data_17;
    assign token_17_36 = token_out_vec_17[32];

    // Process: ProcessingElement_13_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 18, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_18 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_18),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_18),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_18),
        .token_in_vec(token_in_vec_18),
        .dl_detect_in(dl_detect_out),
        .origin(origin[18]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_18),
        .out_chan_dep_data(out_chan_dep_data_18),
        .token_out_vec(token_out_vec_18),
        .dl_detect_out(dl_in_vec[18]));

    assign proc_18_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_12_blk_n) | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_12_blk_n) | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_WriteC_Flattened_fu_179.cPipes_12_blk_n);
    assign proc_18_data_PIPO_blk[0] = 1'b0;
    assign proc_18_start_FIFO_blk[0] = 1'b0;
    assign proc_18_TLF_FIFO_blk[0] = 1'b0;
    assign proc_18_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_18_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_18[0] = dl_detect_out ? proc_dep_vld_vec_18_reg[0] : (proc_18_data_FIFO_blk[0] | proc_18_data_PIPO_blk[0] | proc_18_start_FIFO_blk[0] | proc_18_TLF_FIFO_blk[0] | proc_18_input_sync_blk[0] | proc_18_output_sync_blk[0]);
    assign proc_18_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_13_blk_n) | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_13_blk_n) | (~ProcessingElement_13_U0.grp_ProcessingElement_13_Pipeline_WriteC_Flattened_fu_179.cPipes_13_blk_n);
    assign proc_18_data_PIPO_blk[1] = 1'b0;
    assign proc_18_start_FIFO_blk[1] = 1'b0;
    assign proc_18_TLF_FIFO_blk[1] = 1'b0;
    assign proc_18_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_18_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_18[1] = dl_detect_out ? proc_dep_vld_vec_18_reg[1] : (proc_18_data_FIFO_blk[1] | proc_18_data_PIPO_blk[1] | proc_18_start_FIFO_blk[1] | proc_18_TLF_FIFO_blk[1] | proc_18_input_sync_blk[1] | proc_18_output_sync_blk[1]);
    assign proc_18_data_FIFO_blk[2] = 1'b0;
    assign proc_18_data_PIPO_blk[2] = 1'b0;
    assign proc_18_start_FIFO_blk[2] = 1'b0;
    assign proc_18_TLF_FIFO_blk[2] = 1'b0;
    assign proc_18_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_18_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_18[2] = dl_detect_out ? proc_dep_vld_vec_18_reg[2] : (proc_18_data_FIFO_blk[2] | proc_18_data_PIPO_blk[2] | proc_18_start_FIFO_blk[2] | proc_18_TLF_FIFO_blk[2] | proc_18_input_sync_blk[2] | proc_18_output_sync_blk[2]);
    assign proc_18_data_FIFO_blk[3] = 1'b0;
    assign proc_18_data_PIPO_blk[3] = 1'b0;
    assign proc_18_start_FIFO_blk[3] = 1'b0;
    assign proc_18_TLF_FIFO_blk[3] = 1'b0;
    assign proc_18_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_18_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_18[3] = dl_detect_out ? proc_dep_vld_vec_18_reg[3] : (proc_18_data_FIFO_blk[3] | proc_18_data_PIPO_blk[3] | proc_18_start_FIFO_blk[3] | proc_18_TLF_FIFO_blk[3] | proc_18_input_sync_blk[3] | proc_18_output_sync_blk[3]);
    assign proc_18_data_FIFO_blk[4] = 1'b0;
    assign proc_18_data_PIPO_blk[4] = 1'b0;
    assign proc_18_start_FIFO_blk[4] = 1'b0;
    assign proc_18_TLF_FIFO_blk[4] = 1'b0;
    assign proc_18_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_18_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_18[4] = dl_detect_out ? proc_dep_vld_vec_18_reg[4] : (proc_18_data_FIFO_blk[4] | proc_18_data_PIPO_blk[4] | proc_18_start_FIFO_blk[4] | proc_18_TLF_FIFO_blk[4] | proc_18_input_sync_blk[4] | proc_18_output_sync_blk[4]);
    assign proc_18_data_FIFO_blk[5] = 1'b0;
    assign proc_18_data_PIPO_blk[5] = 1'b0;
    assign proc_18_start_FIFO_blk[5] = 1'b0;
    assign proc_18_TLF_FIFO_blk[5] = 1'b0;
    assign proc_18_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_18_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_18[5] = dl_detect_out ? proc_dep_vld_vec_18_reg[5] : (proc_18_data_FIFO_blk[5] | proc_18_data_PIPO_blk[5] | proc_18_start_FIFO_blk[5] | proc_18_TLF_FIFO_blk[5] | proc_18_input_sync_blk[5] | proc_18_output_sync_blk[5]);
    assign proc_18_data_FIFO_blk[6] = 1'b0;
    assign proc_18_data_PIPO_blk[6] = 1'b0;
    assign proc_18_start_FIFO_blk[6] = 1'b0;
    assign proc_18_TLF_FIFO_blk[6] = 1'b0;
    assign proc_18_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_18_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_18[6] = dl_detect_out ? proc_dep_vld_vec_18_reg[6] : (proc_18_data_FIFO_blk[6] | proc_18_data_PIPO_blk[6] | proc_18_start_FIFO_blk[6] | proc_18_TLF_FIFO_blk[6] | proc_18_input_sync_blk[6] | proc_18_output_sync_blk[6]);
    assign proc_18_data_FIFO_blk[7] = 1'b0;
    assign proc_18_data_PIPO_blk[7] = 1'b0;
    assign proc_18_start_FIFO_blk[7] = 1'b0;
    assign proc_18_TLF_FIFO_blk[7] = 1'b0;
    assign proc_18_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_18_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_18[7] = dl_detect_out ? proc_dep_vld_vec_18_reg[7] : (proc_18_data_FIFO_blk[7] | proc_18_data_PIPO_blk[7] | proc_18_start_FIFO_blk[7] | proc_18_TLF_FIFO_blk[7] | proc_18_input_sync_blk[7] | proc_18_output_sync_blk[7]);
    assign proc_18_data_FIFO_blk[8] = 1'b0;
    assign proc_18_data_PIPO_blk[8] = 1'b0;
    assign proc_18_start_FIFO_blk[8] = 1'b0;
    assign proc_18_TLF_FIFO_blk[8] = 1'b0;
    assign proc_18_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_18_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_18[8] = dl_detect_out ? proc_dep_vld_vec_18_reg[8] : (proc_18_data_FIFO_blk[8] | proc_18_data_PIPO_blk[8] | proc_18_start_FIFO_blk[8] | proc_18_TLF_FIFO_blk[8] | proc_18_input_sync_blk[8] | proc_18_output_sync_blk[8]);
    assign proc_18_data_FIFO_blk[9] = 1'b0;
    assign proc_18_data_PIPO_blk[9] = 1'b0;
    assign proc_18_start_FIFO_blk[9] = 1'b0;
    assign proc_18_TLF_FIFO_blk[9] = 1'b0;
    assign proc_18_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_18_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_18[9] = dl_detect_out ? proc_dep_vld_vec_18_reg[9] : (proc_18_data_FIFO_blk[9] | proc_18_data_PIPO_blk[9] | proc_18_start_FIFO_blk[9] | proc_18_TLF_FIFO_blk[9] | proc_18_input_sync_blk[9] | proc_18_output_sync_blk[9]);
    assign proc_18_data_FIFO_blk[10] = 1'b0;
    assign proc_18_data_PIPO_blk[10] = 1'b0;
    assign proc_18_start_FIFO_blk[10] = 1'b0;
    assign proc_18_TLF_FIFO_blk[10] = 1'b0;
    assign proc_18_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_18_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_18[10] = dl_detect_out ? proc_dep_vld_vec_18_reg[10] : (proc_18_data_FIFO_blk[10] | proc_18_data_PIPO_blk[10] | proc_18_start_FIFO_blk[10] | proc_18_TLF_FIFO_blk[10] | proc_18_input_sync_blk[10] | proc_18_output_sync_blk[10]);
    assign proc_18_data_FIFO_blk[11] = 1'b0;
    assign proc_18_data_PIPO_blk[11] = 1'b0;
    assign proc_18_start_FIFO_blk[11] = 1'b0;
    assign proc_18_TLF_FIFO_blk[11] = 1'b0;
    assign proc_18_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_18_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_18[11] = dl_detect_out ? proc_dep_vld_vec_18_reg[11] : (proc_18_data_FIFO_blk[11] | proc_18_data_PIPO_blk[11] | proc_18_start_FIFO_blk[11] | proc_18_TLF_FIFO_blk[11] | proc_18_input_sync_blk[11] | proc_18_output_sync_blk[11]);
    assign proc_18_data_FIFO_blk[12] = 1'b0;
    assign proc_18_data_PIPO_blk[12] = 1'b0;
    assign proc_18_start_FIFO_blk[12] = 1'b0;
    assign proc_18_TLF_FIFO_blk[12] = 1'b0;
    assign proc_18_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_18_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_18[12] = dl_detect_out ? proc_dep_vld_vec_18_reg[12] : (proc_18_data_FIFO_blk[12] | proc_18_data_PIPO_blk[12] | proc_18_start_FIFO_blk[12] | proc_18_TLF_FIFO_blk[12] | proc_18_input_sync_blk[12] | proc_18_output_sync_blk[12]);
    assign proc_18_data_FIFO_blk[13] = 1'b0;
    assign proc_18_data_PIPO_blk[13] = 1'b0;
    assign proc_18_start_FIFO_blk[13] = 1'b0;
    assign proc_18_TLF_FIFO_blk[13] = 1'b0;
    assign proc_18_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_18_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_18[13] = dl_detect_out ? proc_dep_vld_vec_18_reg[13] : (proc_18_data_FIFO_blk[13] | proc_18_data_PIPO_blk[13] | proc_18_start_FIFO_blk[13] | proc_18_TLF_FIFO_blk[13] | proc_18_input_sync_blk[13] | proc_18_output_sync_blk[13]);
    assign proc_18_data_FIFO_blk[14] = 1'b0;
    assign proc_18_data_PIPO_blk[14] = 1'b0;
    assign proc_18_start_FIFO_blk[14] = 1'b0;
    assign proc_18_TLF_FIFO_blk[14] = 1'b0;
    assign proc_18_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_18_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_18[14] = dl_detect_out ? proc_dep_vld_vec_18_reg[14] : (proc_18_data_FIFO_blk[14] | proc_18_data_PIPO_blk[14] | proc_18_start_FIFO_blk[14] | proc_18_TLF_FIFO_blk[14] | proc_18_input_sync_blk[14] | proc_18_output_sync_blk[14]);
    assign proc_18_data_FIFO_blk[15] = 1'b0;
    assign proc_18_data_PIPO_blk[15] = 1'b0;
    assign proc_18_start_FIFO_blk[15] = 1'b0;
    assign proc_18_TLF_FIFO_blk[15] = 1'b0;
    assign proc_18_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_18_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_18[15] = dl_detect_out ? proc_dep_vld_vec_18_reg[15] : (proc_18_data_FIFO_blk[15] | proc_18_data_PIPO_blk[15] | proc_18_start_FIFO_blk[15] | proc_18_TLF_FIFO_blk[15] | proc_18_input_sync_blk[15] | proc_18_output_sync_blk[15]);
    assign proc_18_data_FIFO_blk[16] = 1'b0;
    assign proc_18_data_PIPO_blk[16] = 1'b0;
    assign proc_18_start_FIFO_blk[16] = 1'b0;
    assign proc_18_TLF_FIFO_blk[16] = 1'b0;
    assign proc_18_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_18_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_18[16] = dl_detect_out ? proc_dep_vld_vec_18_reg[16] : (proc_18_data_FIFO_blk[16] | proc_18_data_PIPO_blk[16] | proc_18_start_FIFO_blk[16] | proc_18_TLF_FIFO_blk[16] | proc_18_input_sync_blk[16] | proc_18_output_sync_blk[16]);
    assign proc_18_data_FIFO_blk[17] = 1'b0;
    assign proc_18_data_PIPO_blk[17] = 1'b0;
    assign proc_18_start_FIFO_blk[17] = 1'b0;
    assign proc_18_TLF_FIFO_blk[17] = 1'b0;
    assign proc_18_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_18_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_18[17] = dl_detect_out ? proc_dep_vld_vec_18_reg[17] : (proc_18_data_FIFO_blk[17] | proc_18_data_PIPO_blk[17] | proc_18_start_FIFO_blk[17] | proc_18_TLF_FIFO_blk[17] | proc_18_input_sync_blk[17] | proc_18_output_sync_blk[17]);
    assign proc_18_data_FIFO_blk[18] = 1'b0;
    assign proc_18_data_PIPO_blk[18] = 1'b0;
    assign proc_18_start_FIFO_blk[18] = 1'b0;
    assign proc_18_TLF_FIFO_blk[18] = 1'b0;
    assign proc_18_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_18_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_18[18] = dl_detect_out ? proc_dep_vld_vec_18_reg[18] : (proc_18_data_FIFO_blk[18] | proc_18_data_PIPO_blk[18] | proc_18_start_FIFO_blk[18] | proc_18_TLF_FIFO_blk[18] | proc_18_input_sync_blk[18] | proc_18_output_sync_blk[18]);
    assign proc_18_data_FIFO_blk[19] = 1'b0;
    assign proc_18_data_PIPO_blk[19] = 1'b0;
    assign proc_18_start_FIFO_blk[19] = 1'b0;
    assign proc_18_TLF_FIFO_blk[19] = 1'b0;
    assign proc_18_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_18_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_18[19] = dl_detect_out ? proc_dep_vld_vec_18_reg[19] : (proc_18_data_FIFO_blk[19] | proc_18_data_PIPO_blk[19] | proc_18_start_FIFO_blk[19] | proc_18_TLF_FIFO_blk[19] | proc_18_input_sync_blk[19] | proc_18_output_sync_blk[19]);
    assign proc_18_data_FIFO_blk[20] = 1'b0;
    assign proc_18_data_PIPO_blk[20] = 1'b0;
    assign proc_18_start_FIFO_blk[20] = 1'b0;
    assign proc_18_TLF_FIFO_blk[20] = 1'b0;
    assign proc_18_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_18_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_18[20] = dl_detect_out ? proc_dep_vld_vec_18_reg[20] : (proc_18_data_FIFO_blk[20] | proc_18_data_PIPO_blk[20] | proc_18_start_FIFO_blk[20] | proc_18_TLF_FIFO_blk[20] | proc_18_input_sync_blk[20] | proc_18_output_sync_blk[20]);
    assign proc_18_data_FIFO_blk[21] = 1'b0;
    assign proc_18_data_PIPO_blk[21] = 1'b0;
    assign proc_18_start_FIFO_blk[21] = 1'b0;
    assign proc_18_TLF_FIFO_blk[21] = 1'b0;
    assign proc_18_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_18_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_18[21] = dl_detect_out ? proc_dep_vld_vec_18_reg[21] : (proc_18_data_FIFO_blk[21] | proc_18_data_PIPO_blk[21] | proc_18_start_FIFO_blk[21] | proc_18_TLF_FIFO_blk[21] | proc_18_input_sync_blk[21] | proc_18_output_sync_blk[21]);
    assign proc_18_data_FIFO_blk[22] = 1'b0;
    assign proc_18_data_PIPO_blk[22] = 1'b0;
    assign proc_18_start_FIFO_blk[22] = 1'b0;
    assign proc_18_TLF_FIFO_blk[22] = 1'b0;
    assign proc_18_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_18_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_18[22] = dl_detect_out ? proc_dep_vld_vec_18_reg[22] : (proc_18_data_FIFO_blk[22] | proc_18_data_PIPO_blk[22] | proc_18_start_FIFO_blk[22] | proc_18_TLF_FIFO_blk[22] | proc_18_input_sync_blk[22] | proc_18_output_sync_blk[22]);
    assign proc_18_data_FIFO_blk[23] = 1'b0;
    assign proc_18_data_PIPO_blk[23] = 1'b0;
    assign proc_18_start_FIFO_blk[23] = 1'b0;
    assign proc_18_TLF_FIFO_blk[23] = 1'b0;
    assign proc_18_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_18_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_18[23] = dl_detect_out ? proc_dep_vld_vec_18_reg[23] : (proc_18_data_FIFO_blk[23] | proc_18_data_PIPO_blk[23] | proc_18_start_FIFO_blk[23] | proc_18_TLF_FIFO_blk[23] | proc_18_input_sync_blk[23] | proc_18_output_sync_blk[23]);
    assign proc_18_data_FIFO_blk[24] = 1'b0;
    assign proc_18_data_PIPO_blk[24] = 1'b0;
    assign proc_18_start_FIFO_blk[24] = 1'b0;
    assign proc_18_TLF_FIFO_blk[24] = 1'b0;
    assign proc_18_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_18_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_18[24] = dl_detect_out ? proc_dep_vld_vec_18_reg[24] : (proc_18_data_FIFO_blk[24] | proc_18_data_PIPO_blk[24] | proc_18_start_FIFO_blk[24] | proc_18_TLF_FIFO_blk[24] | proc_18_input_sync_blk[24] | proc_18_output_sync_blk[24]);
    assign proc_18_data_FIFO_blk[25] = 1'b0;
    assign proc_18_data_PIPO_blk[25] = 1'b0;
    assign proc_18_start_FIFO_blk[25] = 1'b0;
    assign proc_18_TLF_FIFO_blk[25] = 1'b0;
    assign proc_18_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_18_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_18[25] = dl_detect_out ? proc_dep_vld_vec_18_reg[25] : (proc_18_data_FIFO_blk[25] | proc_18_data_PIPO_blk[25] | proc_18_start_FIFO_blk[25] | proc_18_TLF_FIFO_blk[25] | proc_18_input_sync_blk[25] | proc_18_output_sync_blk[25]);
    assign proc_18_data_FIFO_blk[26] = 1'b0;
    assign proc_18_data_PIPO_blk[26] = 1'b0;
    assign proc_18_start_FIFO_blk[26] = 1'b0;
    assign proc_18_TLF_FIFO_blk[26] = 1'b0;
    assign proc_18_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_18_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_18[26] = dl_detect_out ? proc_dep_vld_vec_18_reg[26] : (proc_18_data_FIFO_blk[26] | proc_18_data_PIPO_blk[26] | proc_18_start_FIFO_blk[26] | proc_18_TLF_FIFO_blk[26] | proc_18_input_sync_blk[26] | proc_18_output_sync_blk[26]);
    assign proc_18_data_FIFO_blk[27] = 1'b0;
    assign proc_18_data_PIPO_blk[27] = 1'b0;
    assign proc_18_start_FIFO_blk[27] = 1'b0;
    assign proc_18_TLF_FIFO_blk[27] = 1'b0;
    assign proc_18_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_18_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_18[27] = dl_detect_out ? proc_dep_vld_vec_18_reg[27] : (proc_18_data_FIFO_blk[27] | proc_18_data_PIPO_blk[27] | proc_18_start_FIFO_blk[27] | proc_18_TLF_FIFO_blk[27] | proc_18_input_sync_blk[27] | proc_18_output_sync_blk[27]);
    assign proc_18_data_FIFO_blk[28] = 1'b0;
    assign proc_18_data_PIPO_blk[28] = 1'b0;
    assign proc_18_start_FIFO_blk[28] = 1'b0;
    assign proc_18_TLF_FIFO_blk[28] = 1'b0;
    assign proc_18_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_18_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_18[28] = dl_detect_out ? proc_dep_vld_vec_18_reg[28] : (proc_18_data_FIFO_blk[28] | proc_18_data_PIPO_blk[28] | proc_18_start_FIFO_blk[28] | proc_18_TLF_FIFO_blk[28] | proc_18_input_sync_blk[28] | proc_18_output_sync_blk[28]);
    assign proc_18_data_FIFO_blk[29] = 1'b0;
    assign proc_18_data_PIPO_blk[29] = 1'b0;
    assign proc_18_start_FIFO_blk[29] = 1'b0;
    assign proc_18_TLF_FIFO_blk[29] = 1'b0;
    assign proc_18_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_18_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_18[29] = dl_detect_out ? proc_dep_vld_vec_18_reg[29] : (proc_18_data_FIFO_blk[29] | proc_18_data_PIPO_blk[29] | proc_18_start_FIFO_blk[29] | proc_18_TLF_FIFO_blk[29] | proc_18_input_sync_blk[29] | proc_18_output_sync_blk[29]);
    assign proc_18_data_FIFO_blk[30] = 1'b0;
    assign proc_18_data_PIPO_blk[30] = 1'b0;
    assign proc_18_start_FIFO_blk[30] = 1'b0;
    assign proc_18_TLF_FIFO_blk[30] = 1'b0;
    assign proc_18_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_18_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_18[30] = dl_detect_out ? proc_dep_vld_vec_18_reg[30] : (proc_18_data_FIFO_blk[30] | proc_18_data_PIPO_blk[30] | proc_18_start_FIFO_blk[30] | proc_18_TLF_FIFO_blk[30] | proc_18_input_sync_blk[30] | proc_18_output_sync_blk[30]);
    assign proc_18_data_FIFO_blk[31] = 1'b0;
    assign proc_18_data_PIPO_blk[31] = 1'b0;
    assign proc_18_start_FIFO_blk[31] = 1'b0;
    assign proc_18_TLF_FIFO_blk[31] = 1'b0;
    assign proc_18_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_18_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_18[31] = dl_detect_out ? proc_dep_vld_vec_18_reg[31] : (proc_18_data_FIFO_blk[31] | proc_18_data_PIPO_blk[31] | proc_18_start_FIFO_blk[31] | proc_18_TLF_FIFO_blk[31] | proc_18_input_sync_blk[31] | proc_18_output_sync_blk[31]);
    assign proc_18_data_FIFO_blk[32] = 1'b0;
    assign proc_18_data_PIPO_blk[32] = 1'b0;
    assign proc_18_start_FIFO_blk[32] = 1'b0;
    assign proc_18_TLF_FIFO_blk[32] = 1'b0;
    assign proc_18_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_13_U0_ap_ready & ProcessingElement_13_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_18_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_18[32] = dl_detect_out ? proc_dep_vld_vec_18_reg[32] : (proc_18_data_FIFO_blk[32] | proc_18_data_PIPO_blk[32] | proc_18_start_FIFO_blk[32] | proc_18_TLF_FIFO_blk[32] | proc_18_input_sync_blk[32] | proc_18_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_18_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_18_reg <= proc_dep_vld_vec_18;
        end
    end
    assign in_chan_dep_vld_vec_18[0] = dep_chan_vld_0_18;
    assign in_chan_dep_data_vec_18[39 : 0] = dep_chan_data_0_18;
    assign token_in_vec_18[0] = token_0_18;
    assign in_chan_dep_vld_vec_18[1] = dep_chan_vld_1_18;
    assign in_chan_dep_data_vec_18[79 : 40] = dep_chan_data_1_18;
    assign token_in_vec_18[1] = token_1_18;
    assign in_chan_dep_vld_vec_18[2] = dep_chan_vld_3_18;
    assign in_chan_dep_data_vec_18[119 : 80] = dep_chan_data_3_18;
    assign token_in_vec_18[2] = token_3_18;
    assign in_chan_dep_vld_vec_18[3] = dep_chan_vld_6_18;
    assign in_chan_dep_data_vec_18[159 : 120] = dep_chan_data_6_18;
    assign token_in_vec_18[3] = token_6_18;
    assign in_chan_dep_vld_vec_18[4] = dep_chan_vld_7_18;
    assign in_chan_dep_data_vec_18[199 : 160] = dep_chan_data_7_18;
    assign token_in_vec_18[4] = token_7_18;
    assign in_chan_dep_vld_vec_18[5] = dep_chan_vld_8_18;
    assign in_chan_dep_data_vec_18[239 : 200] = dep_chan_data_8_18;
    assign token_in_vec_18[5] = token_8_18;
    assign in_chan_dep_vld_vec_18[6] = dep_chan_vld_9_18;
    assign in_chan_dep_data_vec_18[279 : 240] = dep_chan_data_9_18;
    assign token_in_vec_18[6] = token_9_18;
    assign in_chan_dep_vld_vec_18[7] = dep_chan_vld_10_18;
    assign in_chan_dep_data_vec_18[319 : 280] = dep_chan_data_10_18;
    assign token_in_vec_18[7] = token_10_18;
    assign in_chan_dep_vld_vec_18[8] = dep_chan_vld_11_18;
    assign in_chan_dep_data_vec_18[359 : 320] = dep_chan_data_11_18;
    assign token_in_vec_18[8] = token_11_18;
    assign in_chan_dep_vld_vec_18[9] = dep_chan_vld_12_18;
    assign in_chan_dep_data_vec_18[399 : 360] = dep_chan_data_12_18;
    assign token_in_vec_18[9] = token_12_18;
    assign in_chan_dep_vld_vec_18[10] = dep_chan_vld_13_18;
    assign in_chan_dep_data_vec_18[439 : 400] = dep_chan_data_13_18;
    assign token_in_vec_18[10] = token_13_18;
    assign in_chan_dep_vld_vec_18[11] = dep_chan_vld_14_18;
    assign in_chan_dep_data_vec_18[479 : 440] = dep_chan_data_14_18;
    assign token_in_vec_18[11] = token_14_18;
    assign in_chan_dep_vld_vec_18[12] = dep_chan_vld_15_18;
    assign in_chan_dep_data_vec_18[519 : 480] = dep_chan_data_15_18;
    assign token_in_vec_18[12] = token_15_18;
    assign in_chan_dep_vld_vec_18[13] = dep_chan_vld_16_18;
    assign in_chan_dep_data_vec_18[559 : 520] = dep_chan_data_16_18;
    assign token_in_vec_18[13] = token_16_18;
    assign in_chan_dep_vld_vec_18[14] = dep_chan_vld_17_18;
    assign in_chan_dep_data_vec_18[599 : 560] = dep_chan_data_17_18;
    assign token_in_vec_18[14] = token_17_18;
    assign in_chan_dep_vld_vec_18[15] = dep_chan_vld_19_18;
    assign in_chan_dep_data_vec_18[639 : 600] = dep_chan_data_19_18;
    assign token_in_vec_18[15] = token_19_18;
    assign in_chan_dep_vld_vec_18[16] = dep_chan_vld_20_18;
    assign in_chan_dep_data_vec_18[679 : 640] = dep_chan_data_20_18;
    assign token_in_vec_18[16] = token_20_18;
    assign in_chan_dep_vld_vec_18[17] = dep_chan_vld_21_18;
    assign in_chan_dep_data_vec_18[719 : 680] = dep_chan_data_21_18;
    assign token_in_vec_18[17] = token_21_18;
    assign in_chan_dep_vld_vec_18[18] = dep_chan_vld_22_18;
    assign in_chan_dep_data_vec_18[759 : 720] = dep_chan_data_22_18;
    assign token_in_vec_18[18] = token_22_18;
    assign in_chan_dep_vld_vec_18[19] = dep_chan_vld_23_18;
    assign in_chan_dep_data_vec_18[799 : 760] = dep_chan_data_23_18;
    assign token_in_vec_18[19] = token_23_18;
    assign in_chan_dep_vld_vec_18[20] = dep_chan_vld_24_18;
    assign in_chan_dep_data_vec_18[839 : 800] = dep_chan_data_24_18;
    assign token_in_vec_18[20] = token_24_18;
    assign in_chan_dep_vld_vec_18[21] = dep_chan_vld_25_18;
    assign in_chan_dep_data_vec_18[879 : 840] = dep_chan_data_25_18;
    assign token_in_vec_18[21] = token_25_18;
    assign in_chan_dep_vld_vec_18[22] = dep_chan_vld_26_18;
    assign in_chan_dep_data_vec_18[919 : 880] = dep_chan_data_26_18;
    assign token_in_vec_18[22] = token_26_18;
    assign in_chan_dep_vld_vec_18[23] = dep_chan_vld_27_18;
    assign in_chan_dep_data_vec_18[959 : 920] = dep_chan_data_27_18;
    assign token_in_vec_18[23] = token_27_18;
    assign in_chan_dep_vld_vec_18[24] = dep_chan_vld_28_18;
    assign in_chan_dep_data_vec_18[999 : 960] = dep_chan_data_28_18;
    assign token_in_vec_18[24] = token_28_18;
    assign in_chan_dep_vld_vec_18[25] = dep_chan_vld_29_18;
    assign in_chan_dep_data_vec_18[1039 : 1000] = dep_chan_data_29_18;
    assign token_in_vec_18[25] = token_29_18;
    assign in_chan_dep_vld_vec_18[26] = dep_chan_vld_30_18;
    assign in_chan_dep_data_vec_18[1079 : 1040] = dep_chan_data_30_18;
    assign token_in_vec_18[26] = token_30_18;
    assign in_chan_dep_vld_vec_18[27] = dep_chan_vld_31_18;
    assign in_chan_dep_data_vec_18[1119 : 1080] = dep_chan_data_31_18;
    assign token_in_vec_18[27] = token_31_18;
    assign in_chan_dep_vld_vec_18[28] = dep_chan_vld_32_18;
    assign in_chan_dep_data_vec_18[1159 : 1120] = dep_chan_data_32_18;
    assign token_in_vec_18[28] = token_32_18;
    assign in_chan_dep_vld_vec_18[29] = dep_chan_vld_33_18;
    assign in_chan_dep_data_vec_18[1199 : 1160] = dep_chan_data_33_18;
    assign token_in_vec_18[29] = token_33_18;
    assign in_chan_dep_vld_vec_18[30] = dep_chan_vld_34_18;
    assign in_chan_dep_data_vec_18[1239 : 1200] = dep_chan_data_34_18;
    assign token_in_vec_18[30] = token_34_18;
    assign in_chan_dep_vld_vec_18[31] = dep_chan_vld_35_18;
    assign in_chan_dep_data_vec_18[1279 : 1240] = dep_chan_data_35_18;
    assign token_in_vec_18[31] = token_35_18;
    assign in_chan_dep_vld_vec_18[32] = dep_chan_vld_36_18;
    assign in_chan_dep_data_vec_18[1319 : 1280] = dep_chan_data_36_18;
    assign token_in_vec_18[32] = token_36_18;
    assign dep_chan_vld_18_17 = out_chan_dep_vld_vec_18[0];
    assign dep_chan_data_18_17 = out_chan_dep_data_18;
    assign token_18_17 = token_out_vec_18[0];
    assign dep_chan_vld_18_19 = out_chan_dep_vld_vec_18[1];
    assign dep_chan_data_18_19 = out_chan_dep_data_18;
    assign token_18_19 = token_out_vec_18[1];
    assign dep_chan_vld_18_0 = out_chan_dep_vld_vec_18[2];
    assign dep_chan_data_18_0 = out_chan_dep_data_18;
    assign token_18_0 = token_out_vec_18[2];
    assign dep_chan_vld_18_1 = out_chan_dep_vld_vec_18[3];
    assign dep_chan_data_18_1 = out_chan_dep_data_18;
    assign token_18_1 = token_out_vec_18[3];
    assign dep_chan_vld_18_3 = out_chan_dep_vld_vec_18[4];
    assign dep_chan_data_18_3 = out_chan_dep_data_18;
    assign token_18_3 = token_out_vec_18[4];
    assign dep_chan_vld_18_6 = out_chan_dep_vld_vec_18[5];
    assign dep_chan_data_18_6 = out_chan_dep_data_18;
    assign token_18_6 = token_out_vec_18[5];
    assign dep_chan_vld_18_7 = out_chan_dep_vld_vec_18[6];
    assign dep_chan_data_18_7 = out_chan_dep_data_18;
    assign token_18_7 = token_out_vec_18[6];
    assign dep_chan_vld_18_8 = out_chan_dep_vld_vec_18[7];
    assign dep_chan_data_18_8 = out_chan_dep_data_18;
    assign token_18_8 = token_out_vec_18[7];
    assign dep_chan_vld_18_9 = out_chan_dep_vld_vec_18[8];
    assign dep_chan_data_18_9 = out_chan_dep_data_18;
    assign token_18_9 = token_out_vec_18[8];
    assign dep_chan_vld_18_10 = out_chan_dep_vld_vec_18[9];
    assign dep_chan_data_18_10 = out_chan_dep_data_18;
    assign token_18_10 = token_out_vec_18[9];
    assign dep_chan_vld_18_11 = out_chan_dep_vld_vec_18[10];
    assign dep_chan_data_18_11 = out_chan_dep_data_18;
    assign token_18_11 = token_out_vec_18[10];
    assign dep_chan_vld_18_12 = out_chan_dep_vld_vec_18[11];
    assign dep_chan_data_18_12 = out_chan_dep_data_18;
    assign token_18_12 = token_out_vec_18[11];
    assign dep_chan_vld_18_13 = out_chan_dep_vld_vec_18[12];
    assign dep_chan_data_18_13 = out_chan_dep_data_18;
    assign token_18_13 = token_out_vec_18[12];
    assign dep_chan_vld_18_14 = out_chan_dep_vld_vec_18[13];
    assign dep_chan_data_18_14 = out_chan_dep_data_18;
    assign token_18_14 = token_out_vec_18[13];
    assign dep_chan_vld_18_15 = out_chan_dep_vld_vec_18[14];
    assign dep_chan_data_18_15 = out_chan_dep_data_18;
    assign token_18_15 = token_out_vec_18[14];
    assign dep_chan_vld_18_16 = out_chan_dep_vld_vec_18[15];
    assign dep_chan_data_18_16 = out_chan_dep_data_18;
    assign token_18_16 = token_out_vec_18[15];
    assign dep_chan_vld_18_20 = out_chan_dep_vld_vec_18[16];
    assign dep_chan_data_18_20 = out_chan_dep_data_18;
    assign token_18_20 = token_out_vec_18[16];
    assign dep_chan_vld_18_21 = out_chan_dep_vld_vec_18[17];
    assign dep_chan_data_18_21 = out_chan_dep_data_18;
    assign token_18_21 = token_out_vec_18[17];
    assign dep_chan_vld_18_22 = out_chan_dep_vld_vec_18[18];
    assign dep_chan_data_18_22 = out_chan_dep_data_18;
    assign token_18_22 = token_out_vec_18[18];
    assign dep_chan_vld_18_23 = out_chan_dep_vld_vec_18[19];
    assign dep_chan_data_18_23 = out_chan_dep_data_18;
    assign token_18_23 = token_out_vec_18[19];
    assign dep_chan_vld_18_24 = out_chan_dep_vld_vec_18[20];
    assign dep_chan_data_18_24 = out_chan_dep_data_18;
    assign token_18_24 = token_out_vec_18[20];
    assign dep_chan_vld_18_25 = out_chan_dep_vld_vec_18[21];
    assign dep_chan_data_18_25 = out_chan_dep_data_18;
    assign token_18_25 = token_out_vec_18[21];
    assign dep_chan_vld_18_26 = out_chan_dep_vld_vec_18[22];
    assign dep_chan_data_18_26 = out_chan_dep_data_18;
    assign token_18_26 = token_out_vec_18[22];
    assign dep_chan_vld_18_27 = out_chan_dep_vld_vec_18[23];
    assign dep_chan_data_18_27 = out_chan_dep_data_18;
    assign token_18_27 = token_out_vec_18[23];
    assign dep_chan_vld_18_28 = out_chan_dep_vld_vec_18[24];
    assign dep_chan_data_18_28 = out_chan_dep_data_18;
    assign token_18_28 = token_out_vec_18[24];
    assign dep_chan_vld_18_29 = out_chan_dep_vld_vec_18[25];
    assign dep_chan_data_18_29 = out_chan_dep_data_18;
    assign token_18_29 = token_out_vec_18[25];
    assign dep_chan_vld_18_30 = out_chan_dep_vld_vec_18[26];
    assign dep_chan_data_18_30 = out_chan_dep_data_18;
    assign token_18_30 = token_out_vec_18[26];
    assign dep_chan_vld_18_31 = out_chan_dep_vld_vec_18[27];
    assign dep_chan_data_18_31 = out_chan_dep_data_18;
    assign token_18_31 = token_out_vec_18[27];
    assign dep_chan_vld_18_32 = out_chan_dep_vld_vec_18[28];
    assign dep_chan_data_18_32 = out_chan_dep_data_18;
    assign token_18_32 = token_out_vec_18[28];
    assign dep_chan_vld_18_33 = out_chan_dep_vld_vec_18[29];
    assign dep_chan_data_18_33 = out_chan_dep_data_18;
    assign token_18_33 = token_out_vec_18[29];
    assign dep_chan_vld_18_34 = out_chan_dep_vld_vec_18[30];
    assign dep_chan_data_18_34 = out_chan_dep_data_18;
    assign token_18_34 = token_out_vec_18[30];
    assign dep_chan_vld_18_35 = out_chan_dep_vld_vec_18[31];
    assign dep_chan_data_18_35 = out_chan_dep_data_18;
    assign token_18_35 = token_out_vec_18[31];
    assign dep_chan_vld_18_36 = out_chan_dep_vld_vec_18[32];
    assign dep_chan_data_18_36 = out_chan_dep_data_18;
    assign token_18_36 = token_out_vec_18[32];

    // Process: ProcessingElement_14_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 19, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_19 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_19),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_19),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_19),
        .token_in_vec(token_in_vec_19),
        .dl_detect_in(dl_detect_out),
        .origin(origin[19]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_19),
        .out_chan_dep_data(out_chan_dep_data_19),
        .token_out_vec(token_out_vec_19),
        .dl_detect_out(dl_in_vec[19]));

    assign proc_19_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_13_blk_n) | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_13_blk_n) | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_WriteC_Flattened_fu_179.cPipes_13_blk_n);
    assign proc_19_data_PIPO_blk[0] = 1'b0;
    assign proc_19_start_FIFO_blk[0] = 1'b0;
    assign proc_19_TLF_FIFO_blk[0] = 1'b0;
    assign proc_19_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_19_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_19[0] = dl_detect_out ? proc_dep_vld_vec_19_reg[0] : (proc_19_data_FIFO_blk[0] | proc_19_data_PIPO_blk[0] | proc_19_start_FIFO_blk[0] | proc_19_TLF_FIFO_blk[0] | proc_19_input_sync_blk[0] | proc_19_output_sync_blk[0]);
    assign proc_19_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_14_blk_n) | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_14_blk_n) | (~ProcessingElement_14_U0.grp_ProcessingElement_14_Pipeline_WriteC_Flattened_fu_179.cPipes_14_blk_n);
    assign proc_19_data_PIPO_blk[1] = 1'b0;
    assign proc_19_start_FIFO_blk[1] = 1'b0;
    assign proc_19_TLF_FIFO_blk[1] = 1'b0;
    assign proc_19_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_19_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_19[1] = dl_detect_out ? proc_dep_vld_vec_19_reg[1] : (proc_19_data_FIFO_blk[1] | proc_19_data_PIPO_blk[1] | proc_19_start_FIFO_blk[1] | proc_19_TLF_FIFO_blk[1] | proc_19_input_sync_blk[1] | proc_19_output_sync_blk[1]);
    assign proc_19_data_FIFO_blk[2] = 1'b0;
    assign proc_19_data_PIPO_blk[2] = 1'b0;
    assign proc_19_start_FIFO_blk[2] = 1'b0;
    assign proc_19_TLF_FIFO_blk[2] = 1'b0;
    assign proc_19_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_19_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_19[2] = dl_detect_out ? proc_dep_vld_vec_19_reg[2] : (proc_19_data_FIFO_blk[2] | proc_19_data_PIPO_blk[2] | proc_19_start_FIFO_blk[2] | proc_19_TLF_FIFO_blk[2] | proc_19_input_sync_blk[2] | proc_19_output_sync_blk[2]);
    assign proc_19_data_FIFO_blk[3] = 1'b0;
    assign proc_19_data_PIPO_blk[3] = 1'b0;
    assign proc_19_start_FIFO_blk[3] = 1'b0;
    assign proc_19_TLF_FIFO_blk[3] = 1'b0;
    assign proc_19_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_19_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_19[3] = dl_detect_out ? proc_dep_vld_vec_19_reg[3] : (proc_19_data_FIFO_blk[3] | proc_19_data_PIPO_blk[3] | proc_19_start_FIFO_blk[3] | proc_19_TLF_FIFO_blk[3] | proc_19_input_sync_blk[3] | proc_19_output_sync_blk[3]);
    assign proc_19_data_FIFO_blk[4] = 1'b0;
    assign proc_19_data_PIPO_blk[4] = 1'b0;
    assign proc_19_start_FIFO_blk[4] = 1'b0;
    assign proc_19_TLF_FIFO_blk[4] = 1'b0;
    assign proc_19_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_19_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_19[4] = dl_detect_out ? proc_dep_vld_vec_19_reg[4] : (proc_19_data_FIFO_blk[4] | proc_19_data_PIPO_blk[4] | proc_19_start_FIFO_blk[4] | proc_19_TLF_FIFO_blk[4] | proc_19_input_sync_blk[4] | proc_19_output_sync_blk[4]);
    assign proc_19_data_FIFO_blk[5] = 1'b0;
    assign proc_19_data_PIPO_blk[5] = 1'b0;
    assign proc_19_start_FIFO_blk[5] = 1'b0;
    assign proc_19_TLF_FIFO_blk[5] = 1'b0;
    assign proc_19_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_19_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_19[5] = dl_detect_out ? proc_dep_vld_vec_19_reg[5] : (proc_19_data_FIFO_blk[5] | proc_19_data_PIPO_blk[5] | proc_19_start_FIFO_blk[5] | proc_19_TLF_FIFO_blk[5] | proc_19_input_sync_blk[5] | proc_19_output_sync_blk[5]);
    assign proc_19_data_FIFO_blk[6] = 1'b0;
    assign proc_19_data_PIPO_blk[6] = 1'b0;
    assign proc_19_start_FIFO_blk[6] = 1'b0;
    assign proc_19_TLF_FIFO_blk[6] = 1'b0;
    assign proc_19_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_19_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_19[6] = dl_detect_out ? proc_dep_vld_vec_19_reg[6] : (proc_19_data_FIFO_blk[6] | proc_19_data_PIPO_blk[6] | proc_19_start_FIFO_blk[6] | proc_19_TLF_FIFO_blk[6] | proc_19_input_sync_blk[6] | proc_19_output_sync_blk[6]);
    assign proc_19_data_FIFO_blk[7] = 1'b0;
    assign proc_19_data_PIPO_blk[7] = 1'b0;
    assign proc_19_start_FIFO_blk[7] = 1'b0;
    assign proc_19_TLF_FIFO_blk[7] = 1'b0;
    assign proc_19_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_19_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_19[7] = dl_detect_out ? proc_dep_vld_vec_19_reg[7] : (proc_19_data_FIFO_blk[7] | proc_19_data_PIPO_blk[7] | proc_19_start_FIFO_blk[7] | proc_19_TLF_FIFO_blk[7] | proc_19_input_sync_blk[7] | proc_19_output_sync_blk[7]);
    assign proc_19_data_FIFO_blk[8] = 1'b0;
    assign proc_19_data_PIPO_blk[8] = 1'b0;
    assign proc_19_start_FIFO_blk[8] = 1'b0;
    assign proc_19_TLF_FIFO_blk[8] = 1'b0;
    assign proc_19_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_19_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_19[8] = dl_detect_out ? proc_dep_vld_vec_19_reg[8] : (proc_19_data_FIFO_blk[8] | proc_19_data_PIPO_blk[8] | proc_19_start_FIFO_blk[8] | proc_19_TLF_FIFO_blk[8] | proc_19_input_sync_blk[8] | proc_19_output_sync_blk[8]);
    assign proc_19_data_FIFO_blk[9] = 1'b0;
    assign proc_19_data_PIPO_blk[9] = 1'b0;
    assign proc_19_start_FIFO_blk[9] = 1'b0;
    assign proc_19_TLF_FIFO_blk[9] = 1'b0;
    assign proc_19_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_19_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_19[9] = dl_detect_out ? proc_dep_vld_vec_19_reg[9] : (proc_19_data_FIFO_blk[9] | proc_19_data_PIPO_blk[9] | proc_19_start_FIFO_blk[9] | proc_19_TLF_FIFO_blk[9] | proc_19_input_sync_blk[9] | proc_19_output_sync_blk[9]);
    assign proc_19_data_FIFO_blk[10] = 1'b0;
    assign proc_19_data_PIPO_blk[10] = 1'b0;
    assign proc_19_start_FIFO_blk[10] = 1'b0;
    assign proc_19_TLF_FIFO_blk[10] = 1'b0;
    assign proc_19_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_19_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_19[10] = dl_detect_out ? proc_dep_vld_vec_19_reg[10] : (proc_19_data_FIFO_blk[10] | proc_19_data_PIPO_blk[10] | proc_19_start_FIFO_blk[10] | proc_19_TLF_FIFO_blk[10] | proc_19_input_sync_blk[10] | proc_19_output_sync_blk[10]);
    assign proc_19_data_FIFO_blk[11] = 1'b0;
    assign proc_19_data_PIPO_blk[11] = 1'b0;
    assign proc_19_start_FIFO_blk[11] = 1'b0;
    assign proc_19_TLF_FIFO_blk[11] = 1'b0;
    assign proc_19_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_19_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_19[11] = dl_detect_out ? proc_dep_vld_vec_19_reg[11] : (proc_19_data_FIFO_blk[11] | proc_19_data_PIPO_blk[11] | proc_19_start_FIFO_blk[11] | proc_19_TLF_FIFO_blk[11] | proc_19_input_sync_blk[11] | proc_19_output_sync_blk[11]);
    assign proc_19_data_FIFO_blk[12] = 1'b0;
    assign proc_19_data_PIPO_blk[12] = 1'b0;
    assign proc_19_start_FIFO_blk[12] = 1'b0;
    assign proc_19_TLF_FIFO_blk[12] = 1'b0;
    assign proc_19_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_19_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_19[12] = dl_detect_out ? proc_dep_vld_vec_19_reg[12] : (proc_19_data_FIFO_blk[12] | proc_19_data_PIPO_blk[12] | proc_19_start_FIFO_blk[12] | proc_19_TLF_FIFO_blk[12] | proc_19_input_sync_blk[12] | proc_19_output_sync_blk[12]);
    assign proc_19_data_FIFO_blk[13] = 1'b0;
    assign proc_19_data_PIPO_blk[13] = 1'b0;
    assign proc_19_start_FIFO_blk[13] = 1'b0;
    assign proc_19_TLF_FIFO_blk[13] = 1'b0;
    assign proc_19_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_19_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_19[13] = dl_detect_out ? proc_dep_vld_vec_19_reg[13] : (proc_19_data_FIFO_blk[13] | proc_19_data_PIPO_blk[13] | proc_19_start_FIFO_blk[13] | proc_19_TLF_FIFO_blk[13] | proc_19_input_sync_blk[13] | proc_19_output_sync_blk[13]);
    assign proc_19_data_FIFO_blk[14] = 1'b0;
    assign proc_19_data_PIPO_blk[14] = 1'b0;
    assign proc_19_start_FIFO_blk[14] = 1'b0;
    assign proc_19_TLF_FIFO_blk[14] = 1'b0;
    assign proc_19_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_19_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_19[14] = dl_detect_out ? proc_dep_vld_vec_19_reg[14] : (proc_19_data_FIFO_blk[14] | proc_19_data_PIPO_blk[14] | proc_19_start_FIFO_blk[14] | proc_19_TLF_FIFO_blk[14] | proc_19_input_sync_blk[14] | proc_19_output_sync_blk[14]);
    assign proc_19_data_FIFO_blk[15] = 1'b0;
    assign proc_19_data_PIPO_blk[15] = 1'b0;
    assign proc_19_start_FIFO_blk[15] = 1'b0;
    assign proc_19_TLF_FIFO_blk[15] = 1'b0;
    assign proc_19_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_19_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_19[15] = dl_detect_out ? proc_dep_vld_vec_19_reg[15] : (proc_19_data_FIFO_blk[15] | proc_19_data_PIPO_blk[15] | proc_19_start_FIFO_blk[15] | proc_19_TLF_FIFO_blk[15] | proc_19_input_sync_blk[15] | proc_19_output_sync_blk[15]);
    assign proc_19_data_FIFO_blk[16] = 1'b0;
    assign proc_19_data_PIPO_blk[16] = 1'b0;
    assign proc_19_start_FIFO_blk[16] = 1'b0;
    assign proc_19_TLF_FIFO_blk[16] = 1'b0;
    assign proc_19_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_19_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_19[16] = dl_detect_out ? proc_dep_vld_vec_19_reg[16] : (proc_19_data_FIFO_blk[16] | proc_19_data_PIPO_blk[16] | proc_19_start_FIFO_blk[16] | proc_19_TLF_FIFO_blk[16] | proc_19_input_sync_blk[16] | proc_19_output_sync_blk[16]);
    assign proc_19_data_FIFO_blk[17] = 1'b0;
    assign proc_19_data_PIPO_blk[17] = 1'b0;
    assign proc_19_start_FIFO_blk[17] = 1'b0;
    assign proc_19_TLF_FIFO_blk[17] = 1'b0;
    assign proc_19_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_19_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_19[17] = dl_detect_out ? proc_dep_vld_vec_19_reg[17] : (proc_19_data_FIFO_blk[17] | proc_19_data_PIPO_blk[17] | proc_19_start_FIFO_blk[17] | proc_19_TLF_FIFO_blk[17] | proc_19_input_sync_blk[17] | proc_19_output_sync_blk[17]);
    assign proc_19_data_FIFO_blk[18] = 1'b0;
    assign proc_19_data_PIPO_blk[18] = 1'b0;
    assign proc_19_start_FIFO_blk[18] = 1'b0;
    assign proc_19_TLF_FIFO_blk[18] = 1'b0;
    assign proc_19_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_19_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_19[18] = dl_detect_out ? proc_dep_vld_vec_19_reg[18] : (proc_19_data_FIFO_blk[18] | proc_19_data_PIPO_blk[18] | proc_19_start_FIFO_blk[18] | proc_19_TLF_FIFO_blk[18] | proc_19_input_sync_blk[18] | proc_19_output_sync_blk[18]);
    assign proc_19_data_FIFO_blk[19] = 1'b0;
    assign proc_19_data_PIPO_blk[19] = 1'b0;
    assign proc_19_start_FIFO_blk[19] = 1'b0;
    assign proc_19_TLF_FIFO_blk[19] = 1'b0;
    assign proc_19_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_19_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_19[19] = dl_detect_out ? proc_dep_vld_vec_19_reg[19] : (proc_19_data_FIFO_blk[19] | proc_19_data_PIPO_blk[19] | proc_19_start_FIFO_blk[19] | proc_19_TLF_FIFO_blk[19] | proc_19_input_sync_blk[19] | proc_19_output_sync_blk[19]);
    assign proc_19_data_FIFO_blk[20] = 1'b0;
    assign proc_19_data_PIPO_blk[20] = 1'b0;
    assign proc_19_start_FIFO_blk[20] = 1'b0;
    assign proc_19_TLF_FIFO_blk[20] = 1'b0;
    assign proc_19_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_19_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_19[20] = dl_detect_out ? proc_dep_vld_vec_19_reg[20] : (proc_19_data_FIFO_blk[20] | proc_19_data_PIPO_blk[20] | proc_19_start_FIFO_blk[20] | proc_19_TLF_FIFO_blk[20] | proc_19_input_sync_blk[20] | proc_19_output_sync_blk[20]);
    assign proc_19_data_FIFO_blk[21] = 1'b0;
    assign proc_19_data_PIPO_blk[21] = 1'b0;
    assign proc_19_start_FIFO_blk[21] = 1'b0;
    assign proc_19_TLF_FIFO_blk[21] = 1'b0;
    assign proc_19_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_19_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_19[21] = dl_detect_out ? proc_dep_vld_vec_19_reg[21] : (proc_19_data_FIFO_blk[21] | proc_19_data_PIPO_blk[21] | proc_19_start_FIFO_blk[21] | proc_19_TLF_FIFO_blk[21] | proc_19_input_sync_blk[21] | proc_19_output_sync_blk[21]);
    assign proc_19_data_FIFO_blk[22] = 1'b0;
    assign proc_19_data_PIPO_blk[22] = 1'b0;
    assign proc_19_start_FIFO_blk[22] = 1'b0;
    assign proc_19_TLF_FIFO_blk[22] = 1'b0;
    assign proc_19_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_19_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_19[22] = dl_detect_out ? proc_dep_vld_vec_19_reg[22] : (proc_19_data_FIFO_blk[22] | proc_19_data_PIPO_blk[22] | proc_19_start_FIFO_blk[22] | proc_19_TLF_FIFO_blk[22] | proc_19_input_sync_blk[22] | proc_19_output_sync_blk[22]);
    assign proc_19_data_FIFO_blk[23] = 1'b0;
    assign proc_19_data_PIPO_blk[23] = 1'b0;
    assign proc_19_start_FIFO_blk[23] = 1'b0;
    assign proc_19_TLF_FIFO_blk[23] = 1'b0;
    assign proc_19_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_19_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_19[23] = dl_detect_out ? proc_dep_vld_vec_19_reg[23] : (proc_19_data_FIFO_blk[23] | proc_19_data_PIPO_blk[23] | proc_19_start_FIFO_blk[23] | proc_19_TLF_FIFO_blk[23] | proc_19_input_sync_blk[23] | proc_19_output_sync_blk[23]);
    assign proc_19_data_FIFO_blk[24] = 1'b0;
    assign proc_19_data_PIPO_blk[24] = 1'b0;
    assign proc_19_start_FIFO_blk[24] = 1'b0;
    assign proc_19_TLF_FIFO_blk[24] = 1'b0;
    assign proc_19_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_19_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_19[24] = dl_detect_out ? proc_dep_vld_vec_19_reg[24] : (proc_19_data_FIFO_blk[24] | proc_19_data_PIPO_blk[24] | proc_19_start_FIFO_blk[24] | proc_19_TLF_FIFO_blk[24] | proc_19_input_sync_blk[24] | proc_19_output_sync_blk[24]);
    assign proc_19_data_FIFO_blk[25] = 1'b0;
    assign proc_19_data_PIPO_blk[25] = 1'b0;
    assign proc_19_start_FIFO_blk[25] = 1'b0;
    assign proc_19_TLF_FIFO_blk[25] = 1'b0;
    assign proc_19_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_19_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_19[25] = dl_detect_out ? proc_dep_vld_vec_19_reg[25] : (proc_19_data_FIFO_blk[25] | proc_19_data_PIPO_blk[25] | proc_19_start_FIFO_blk[25] | proc_19_TLF_FIFO_blk[25] | proc_19_input_sync_blk[25] | proc_19_output_sync_blk[25]);
    assign proc_19_data_FIFO_blk[26] = 1'b0;
    assign proc_19_data_PIPO_blk[26] = 1'b0;
    assign proc_19_start_FIFO_blk[26] = 1'b0;
    assign proc_19_TLF_FIFO_blk[26] = 1'b0;
    assign proc_19_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_19_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_19[26] = dl_detect_out ? proc_dep_vld_vec_19_reg[26] : (proc_19_data_FIFO_blk[26] | proc_19_data_PIPO_blk[26] | proc_19_start_FIFO_blk[26] | proc_19_TLF_FIFO_blk[26] | proc_19_input_sync_blk[26] | proc_19_output_sync_blk[26]);
    assign proc_19_data_FIFO_blk[27] = 1'b0;
    assign proc_19_data_PIPO_blk[27] = 1'b0;
    assign proc_19_start_FIFO_blk[27] = 1'b0;
    assign proc_19_TLF_FIFO_blk[27] = 1'b0;
    assign proc_19_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_19_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_19[27] = dl_detect_out ? proc_dep_vld_vec_19_reg[27] : (proc_19_data_FIFO_blk[27] | proc_19_data_PIPO_blk[27] | proc_19_start_FIFO_blk[27] | proc_19_TLF_FIFO_blk[27] | proc_19_input_sync_blk[27] | proc_19_output_sync_blk[27]);
    assign proc_19_data_FIFO_blk[28] = 1'b0;
    assign proc_19_data_PIPO_blk[28] = 1'b0;
    assign proc_19_start_FIFO_blk[28] = 1'b0;
    assign proc_19_TLF_FIFO_blk[28] = 1'b0;
    assign proc_19_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_19_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_19[28] = dl_detect_out ? proc_dep_vld_vec_19_reg[28] : (proc_19_data_FIFO_blk[28] | proc_19_data_PIPO_blk[28] | proc_19_start_FIFO_blk[28] | proc_19_TLF_FIFO_blk[28] | proc_19_input_sync_blk[28] | proc_19_output_sync_blk[28]);
    assign proc_19_data_FIFO_blk[29] = 1'b0;
    assign proc_19_data_PIPO_blk[29] = 1'b0;
    assign proc_19_start_FIFO_blk[29] = 1'b0;
    assign proc_19_TLF_FIFO_blk[29] = 1'b0;
    assign proc_19_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_19_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_19[29] = dl_detect_out ? proc_dep_vld_vec_19_reg[29] : (proc_19_data_FIFO_blk[29] | proc_19_data_PIPO_blk[29] | proc_19_start_FIFO_blk[29] | proc_19_TLF_FIFO_blk[29] | proc_19_input_sync_blk[29] | proc_19_output_sync_blk[29]);
    assign proc_19_data_FIFO_blk[30] = 1'b0;
    assign proc_19_data_PIPO_blk[30] = 1'b0;
    assign proc_19_start_FIFO_blk[30] = 1'b0;
    assign proc_19_TLF_FIFO_blk[30] = 1'b0;
    assign proc_19_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_19_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_19[30] = dl_detect_out ? proc_dep_vld_vec_19_reg[30] : (proc_19_data_FIFO_blk[30] | proc_19_data_PIPO_blk[30] | proc_19_start_FIFO_blk[30] | proc_19_TLF_FIFO_blk[30] | proc_19_input_sync_blk[30] | proc_19_output_sync_blk[30]);
    assign proc_19_data_FIFO_blk[31] = 1'b0;
    assign proc_19_data_PIPO_blk[31] = 1'b0;
    assign proc_19_start_FIFO_blk[31] = 1'b0;
    assign proc_19_TLF_FIFO_blk[31] = 1'b0;
    assign proc_19_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_19_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_19[31] = dl_detect_out ? proc_dep_vld_vec_19_reg[31] : (proc_19_data_FIFO_blk[31] | proc_19_data_PIPO_blk[31] | proc_19_start_FIFO_blk[31] | proc_19_TLF_FIFO_blk[31] | proc_19_input_sync_blk[31] | proc_19_output_sync_blk[31]);
    assign proc_19_data_FIFO_blk[32] = 1'b0;
    assign proc_19_data_PIPO_blk[32] = 1'b0;
    assign proc_19_start_FIFO_blk[32] = 1'b0;
    assign proc_19_TLF_FIFO_blk[32] = 1'b0;
    assign proc_19_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_14_U0_ap_ready & ProcessingElement_14_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_19_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_19[32] = dl_detect_out ? proc_dep_vld_vec_19_reg[32] : (proc_19_data_FIFO_blk[32] | proc_19_data_PIPO_blk[32] | proc_19_start_FIFO_blk[32] | proc_19_TLF_FIFO_blk[32] | proc_19_input_sync_blk[32] | proc_19_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_19_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_19_reg <= proc_dep_vld_vec_19;
        end
    end
    assign in_chan_dep_vld_vec_19[0] = dep_chan_vld_0_19;
    assign in_chan_dep_data_vec_19[39 : 0] = dep_chan_data_0_19;
    assign token_in_vec_19[0] = token_0_19;
    assign in_chan_dep_vld_vec_19[1] = dep_chan_vld_1_19;
    assign in_chan_dep_data_vec_19[79 : 40] = dep_chan_data_1_19;
    assign token_in_vec_19[1] = token_1_19;
    assign in_chan_dep_vld_vec_19[2] = dep_chan_vld_3_19;
    assign in_chan_dep_data_vec_19[119 : 80] = dep_chan_data_3_19;
    assign token_in_vec_19[2] = token_3_19;
    assign in_chan_dep_vld_vec_19[3] = dep_chan_vld_6_19;
    assign in_chan_dep_data_vec_19[159 : 120] = dep_chan_data_6_19;
    assign token_in_vec_19[3] = token_6_19;
    assign in_chan_dep_vld_vec_19[4] = dep_chan_vld_7_19;
    assign in_chan_dep_data_vec_19[199 : 160] = dep_chan_data_7_19;
    assign token_in_vec_19[4] = token_7_19;
    assign in_chan_dep_vld_vec_19[5] = dep_chan_vld_8_19;
    assign in_chan_dep_data_vec_19[239 : 200] = dep_chan_data_8_19;
    assign token_in_vec_19[5] = token_8_19;
    assign in_chan_dep_vld_vec_19[6] = dep_chan_vld_9_19;
    assign in_chan_dep_data_vec_19[279 : 240] = dep_chan_data_9_19;
    assign token_in_vec_19[6] = token_9_19;
    assign in_chan_dep_vld_vec_19[7] = dep_chan_vld_10_19;
    assign in_chan_dep_data_vec_19[319 : 280] = dep_chan_data_10_19;
    assign token_in_vec_19[7] = token_10_19;
    assign in_chan_dep_vld_vec_19[8] = dep_chan_vld_11_19;
    assign in_chan_dep_data_vec_19[359 : 320] = dep_chan_data_11_19;
    assign token_in_vec_19[8] = token_11_19;
    assign in_chan_dep_vld_vec_19[9] = dep_chan_vld_12_19;
    assign in_chan_dep_data_vec_19[399 : 360] = dep_chan_data_12_19;
    assign token_in_vec_19[9] = token_12_19;
    assign in_chan_dep_vld_vec_19[10] = dep_chan_vld_13_19;
    assign in_chan_dep_data_vec_19[439 : 400] = dep_chan_data_13_19;
    assign token_in_vec_19[10] = token_13_19;
    assign in_chan_dep_vld_vec_19[11] = dep_chan_vld_14_19;
    assign in_chan_dep_data_vec_19[479 : 440] = dep_chan_data_14_19;
    assign token_in_vec_19[11] = token_14_19;
    assign in_chan_dep_vld_vec_19[12] = dep_chan_vld_15_19;
    assign in_chan_dep_data_vec_19[519 : 480] = dep_chan_data_15_19;
    assign token_in_vec_19[12] = token_15_19;
    assign in_chan_dep_vld_vec_19[13] = dep_chan_vld_16_19;
    assign in_chan_dep_data_vec_19[559 : 520] = dep_chan_data_16_19;
    assign token_in_vec_19[13] = token_16_19;
    assign in_chan_dep_vld_vec_19[14] = dep_chan_vld_17_19;
    assign in_chan_dep_data_vec_19[599 : 560] = dep_chan_data_17_19;
    assign token_in_vec_19[14] = token_17_19;
    assign in_chan_dep_vld_vec_19[15] = dep_chan_vld_18_19;
    assign in_chan_dep_data_vec_19[639 : 600] = dep_chan_data_18_19;
    assign token_in_vec_19[15] = token_18_19;
    assign in_chan_dep_vld_vec_19[16] = dep_chan_vld_20_19;
    assign in_chan_dep_data_vec_19[679 : 640] = dep_chan_data_20_19;
    assign token_in_vec_19[16] = token_20_19;
    assign in_chan_dep_vld_vec_19[17] = dep_chan_vld_21_19;
    assign in_chan_dep_data_vec_19[719 : 680] = dep_chan_data_21_19;
    assign token_in_vec_19[17] = token_21_19;
    assign in_chan_dep_vld_vec_19[18] = dep_chan_vld_22_19;
    assign in_chan_dep_data_vec_19[759 : 720] = dep_chan_data_22_19;
    assign token_in_vec_19[18] = token_22_19;
    assign in_chan_dep_vld_vec_19[19] = dep_chan_vld_23_19;
    assign in_chan_dep_data_vec_19[799 : 760] = dep_chan_data_23_19;
    assign token_in_vec_19[19] = token_23_19;
    assign in_chan_dep_vld_vec_19[20] = dep_chan_vld_24_19;
    assign in_chan_dep_data_vec_19[839 : 800] = dep_chan_data_24_19;
    assign token_in_vec_19[20] = token_24_19;
    assign in_chan_dep_vld_vec_19[21] = dep_chan_vld_25_19;
    assign in_chan_dep_data_vec_19[879 : 840] = dep_chan_data_25_19;
    assign token_in_vec_19[21] = token_25_19;
    assign in_chan_dep_vld_vec_19[22] = dep_chan_vld_26_19;
    assign in_chan_dep_data_vec_19[919 : 880] = dep_chan_data_26_19;
    assign token_in_vec_19[22] = token_26_19;
    assign in_chan_dep_vld_vec_19[23] = dep_chan_vld_27_19;
    assign in_chan_dep_data_vec_19[959 : 920] = dep_chan_data_27_19;
    assign token_in_vec_19[23] = token_27_19;
    assign in_chan_dep_vld_vec_19[24] = dep_chan_vld_28_19;
    assign in_chan_dep_data_vec_19[999 : 960] = dep_chan_data_28_19;
    assign token_in_vec_19[24] = token_28_19;
    assign in_chan_dep_vld_vec_19[25] = dep_chan_vld_29_19;
    assign in_chan_dep_data_vec_19[1039 : 1000] = dep_chan_data_29_19;
    assign token_in_vec_19[25] = token_29_19;
    assign in_chan_dep_vld_vec_19[26] = dep_chan_vld_30_19;
    assign in_chan_dep_data_vec_19[1079 : 1040] = dep_chan_data_30_19;
    assign token_in_vec_19[26] = token_30_19;
    assign in_chan_dep_vld_vec_19[27] = dep_chan_vld_31_19;
    assign in_chan_dep_data_vec_19[1119 : 1080] = dep_chan_data_31_19;
    assign token_in_vec_19[27] = token_31_19;
    assign in_chan_dep_vld_vec_19[28] = dep_chan_vld_32_19;
    assign in_chan_dep_data_vec_19[1159 : 1120] = dep_chan_data_32_19;
    assign token_in_vec_19[28] = token_32_19;
    assign in_chan_dep_vld_vec_19[29] = dep_chan_vld_33_19;
    assign in_chan_dep_data_vec_19[1199 : 1160] = dep_chan_data_33_19;
    assign token_in_vec_19[29] = token_33_19;
    assign in_chan_dep_vld_vec_19[30] = dep_chan_vld_34_19;
    assign in_chan_dep_data_vec_19[1239 : 1200] = dep_chan_data_34_19;
    assign token_in_vec_19[30] = token_34_19;
    assign in_chan_dep_vld_vec_19[31] = dep_chan_vld_35_19;
    assign in_chan_dep_data_vec_19[1279 : 1240] = dep_chan_data_35_19;
    assign token_in_vec_19[31] = token_35_19;
    assign in_chan_dep_vld_vec_19[32] = dep_chan_vld_36_19;
    assign in_chan_dep_data_vec_19[1319 : 1280] = dep_chan_data_36_19;
    assign token_in_vec_19[32] = token_36_19;
    assign dep_chan_vld_19_18 = out_chan_dep_vld_vec_19[0];
    assign dep_chan_data_19_18 = out_chan_dep_data_19;
    assign token_19_18 = token_out_vec_19[0];
    assign dep_chan_vld_19_20 = out_chan_dep_vld_vec_19[1];
    assign dep_chan_data_19_20 = out_chan_dep_data_19;
    assign token_19_20 = token_out_vec_19[1];
    assign dep_chan_vld_19_0 = out_chan_dep_vld_vec_19[2];
    assign dep_chan_data_19_0 = out_chan_dep_data_19;
    assign token_19_0 = token_out_vec_19[2];
    assign dep_chan_vld_19_1 = out_chan_dep_vld_vec_19[3];
    assign dep_chan_data_19_1 = out_chan_dep_data_19;
    assign token_19_1 = token_out_vec_19[3];
    assign dep_chan_vld_19_3 = out_chan_dep_vld_vec_19[4];
    assign dep_chan_data_19_3 = out_chan_dep_data_19;
    assign token_19_3 = token_out_vec_19[4];
    assign dep_chan_vld_19_6 = out_chan_dep_vld_vec_19[5];
    assign dep_chan_data_19_6 = out_chan_dep_data_19;
    assign token_19_6 = token_out_vec_19[5];
    assign dep_chan_vld_19_7 = out_chan_dep_vld_vec_19[6];
    assign dep_chan_data_19_7 = out_chan_dep_data_19;
    assign token_19_7 = token_out_vec_19[6];
    assign dep_chan_vld_19_8 = out_chan_dep_vld_vec_19[7];
    assign dep_chan_data_19_8 = out_chan_dep_data_19;
    assign token_19_8 = token_out_vec_19[7];
    assign dep_chan_vld_19_9 = out_chan_dep_vld_vec_19[8];
    assign dep_chan_data_19_9 = out_chan_dep_data_19;
    assign token_19_9 = token_out_vec_19[8];
    assign dep_chan_vld_19_10 = out_chan_dep_vld_vec_19[9];
    assign dep_chan_data_19_10 = out_chan_dep_data_19;
    assign token_19_10 = token_out_vec_19[9];
    assign dep_chan_vld_19_11 = out_chan_dep_vld_vec_19[10];
    assign dep_chan_data_19_11 = out_chan_dep_data_19;
    assign token_19_11 = token_out_vec_19[10];
    assign dep_chan_vld_19_12 = out_chan_dep_vld_vec_19[11];
    assign dep_chan_data_19_12 = out_chan_dep_data_19;
    assign token_19_12 = token_out_vec_19[11];
    assign dep_chan_vld_19_13 = out_chan_dep_vld_vec_19[12];
    assign dep_chan_data_19_13 = out_chan_dep_data_19;
    assign token_19_13 = token_out_vec_19[12];
    assign dep_chan_vld_19_14 = out_chan_dep_vld_vec_19[13];
    assign dep_chan_data_19_14 = out_chan_dep_data_19;
    assign token_19_14 = token_out_vec_19[13];
    assign dep_chan_vld_19_15 = out_chan_dep_vld_vec_19[14];
    assign dep_chan_data_19_15 = out_chan_dep_data_19;
    assign token_19_15 = token_out_vec_19[14];
    assign dep_chan_vld_19_16 = out_chan_dep_vld_vec_19[15];
    assign dep_chan_data_19_16 = out_chan_dep_data_19;
    assign token_19_16 = token_out_vec_19[15];
    assign dep_chan_vld_19_17 = out_chan_dep_vld_vec_19[16];
    assign dep_chan_data_19_17 = out_chan_dep_data_19;
    assign token_19_17 = token_out_vec_19[16];
    assign dep_chan_vld_19_21 = out_chan_dep_vld_vec_19[17];
    assign dep_chan_data_19_21 = out_chan_dep_data_19;
    assign token_19_21 = token_out_vec_19[17];
    assign dep_chan_vld_19_22 = out_chan_dep_vld_vec_19[18];
    assign dep_chan_data_19_22 = out_chan_dep_data_19;
    assign token_19_22 = token_out_vec_19[18];
    assign dep_chan_vld_19_23 = out_chan_dep_vld_vec_19[19];
    assign dep_chan_data_19_23 = out_chan_dep_data_19;
    assign token_19_23 = token_out_vec_19[19];
    assign dep_chan_vld_19_24 = out_chan_dep_vld_vec_19[20];
    assign dep_chan_data_19_24 = out_chan_dep_data_19;
    assign token_19_24 = token_out_vec_19[20];
    assign dep_chan_vld_19_25 = out_chan_dep_vld_vec_19[21];
    assign dep_chan_data_19_25 = out_chan_dep_data_19;
    assign token_19_25 = token_out_vec_19[21];
    assign dep_chan_vld_19_26 = out_chan_dep_vld_vec_19[22];
    assign dep_chan_data_19_26 = out_chan_dep_data_19;
    assign token_19_26 = token_out_vec_19[22];
    assign dep_chan_vld_19_27 = out_chan_dep_vld_vec_19[23];
    assign dep_chan_data_19_27 = out_chan_dep_data_19;
    assign token_19_27 = token_out_vec_19[23];
    assign dep_chan_vld_19_28 = out_chan_dep_vld_vec_19[24];
    assign dep_chan_data_19_28 = out_chan_dep_data_19;
    assign token_19_28 = token_out_vec_19[24];
    assign dep_chan_vld_19_29 = out_chan_dep_vld_vec_19[25];
    assign dep_chan_data_19_29 = out_chan_dep_data_19;
    assign token_19_29 = token_out_vec_19[25];
    assign dep_chan_vld_19_30 = out_chan_dep_vld_vec_19[26];
    assign dep_chan_data_19_30 = out_chan_dep_data_19;
    assign token_19_30 = token_out_vec_19[26];
    assign dep_chan_vld_19_31 = out_chan_dep_vld_vec_19[27];
    assign dep_chan_data_19_31 = out_chan_dep_data_19;
    assign token_19_31 = token_out_vec_19[27];
    assign dep_chan_vld_19_32 = out_chan_dep_vld_vec_19[28];
    assign dep_chan_data_19_32 = out_chan_dep_data_19;
    assign token_19_32 = token_out_vec_19[28];
    assign dep_chan_vld_19_33 = out_chan_dep_vld_vec_19[29];
    assign dep_chan_data_19_33 = out_chan_dep_data_19;
    assign token_19_33 = token_out_vec_19[29];
    assign dep_chan_vld_19_34 = out_chan_dep_vld_vec_19[30];
    assign dep_chan_data_19_34 = out_chan_dep_data_19;
    assign token_19_34 = token_out_vec_19[30];
    assign dep_chan_vld_19_35 = out_chan_dep_vld_vec_19[31];
    assign dep_chan_data_19_35 = out_chan_dep_data_19;
    assign token_19_35 = token_out_vec_19[31];
    assign dep_chan_vld_19_36 = out_chan_dep_vld_vec_19[32];
    assign dep_chan_data_19_36 = out_chan_dep_data_19;
    assign token_19_36 = token_out_vec_19[32];

    // Process: ProcessingElement_15_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 20, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_20 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_20),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_20),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_20),
        .token_in_vec(token_in_vec_20),
        .dl_detect_in(dl_detect_out),
        .origin(origin[20]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_20),
        .out_chan_dep_data(out_chan_dep_data_20),
        .token_out_vec(token_out_vec_20),
        .dl_detect_out(dl_in_vec[20]));

    assign proc_20_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_14_blk_n) | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_14_blk_n) | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_WriteC_Flattened_fu_179.cPipes_14_blk_n);
    assign proc_20_data_PIPO_blk[0] = 1'b0;
    assign proc_20_start_FIFO_blk[0] = 1'b0;
    assign proc_20_TLF_FIFO_blk[0] = 1'b0;
    assign proc_20_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_20_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_20[0] = dl_detect_out ? proc_dep_vld_vec_20_reg[0] : (proc_20_data_FIFO_blk[0] | proc_20_data_PIPO_blk[0] | proc_20_start_FIFO_blk[0] | proc_20_TLF_FIFO_blk[0] | proc_20_input_sync_blk[0] | proc_20_output_sync_blk[0]);
    assign proc_20_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_15_blk_n) | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_15_blk_n) | (~ProcessingElement_15_U0.grp_ProcessingElement_15_Pipeline_WriteC_Flattened_fu_179.cPipes_15_blk_n);
    assign proc_20_data_PIPO_blk[1] = 1'b0;
    assign proc_20_start_FIFO_blk[1] = 1'b0;
    assign proc_20_TLF_FIFO_blk[1] = 1'b0;
    assign proc_20_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_20_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_20[1] = dl_detect_out ? proc_dep_vld_vec_20_reg[1] : (proc_20_data_FIFO_blk[1] | proc_20_data_PIPO_blk[1] | proc_20_start_FIFO_blk[1] | proc_20_TLF_FIFO_blk[1] | proc_20_input_sync_blk[1] | proc_20_output_sync_blk[1]);
    assign proc_20_data_FIFO_blk[2] = 1'b0;
    assign proc_20_data_PIPO_blk[2] = 1'b0;
    assign proc_20_start_FIFO_blk[2] = 1'b0;
    assign proc_20_TLF_FIFO_blk[2] = 1'b0;
    assign proc_20_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_20_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_20[2] = dl_detect_out ? proc_dep_vld_vec_20_reg[2] : (proc_20_data_FIFO_blk[2] | proc_20_data_PIPO_blk[2] | proc_20_start_FIFO_blk[2] | proc_20_TLF_FIFO_blk[2] | proc_20_input_sync_blk[2] | proc_20_output_sync_blk[2]);
    assign proc_20_data_FIFO_blk[3] = 1'b0;
    assign proc_20_data_PIPO_blk[3] = 1'b0;
    assign proc_20_start_FIFO_blk[3] = 1'b0;
    assign proc_20_TLF_FIFO_blk[3] = 1'b0;
    assign proc_20_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_20_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_20[3] = dl_detect_out ? proc_dep_vld_vec_20_reg[3] : (proc_20_data_FIFO_blk[3] | proc_20_data_PIPO_blk[3] | proc_20_start_FIFO_blk[3] | proc_20_TLF_FIFO_blk[3] | proc_20_input_sync_blk[3] | proc_20_output_sync_blk[3]);
    assign proc_20_data_FIFO_blk[4] = 1'b0;
    assign proc_20_data_PIPO_blk[4] = 1'b0;
    assign proc_20_start_FIFO_blk[4] = 1'b0;
    assign proc_20_TLF_FIFO_blk[4] = 1'b0;
    assign proc_20_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_20_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_20[4] = dl_detect_out ? proc_dep_vld_vec_20_reg[4] : (proc_20_data_FIFO_blk[4] | proc_20_data_PIPO_blk[4] | proc_20_start_FIFO_blk[4] | proc_20_TLF_FIFO_blk[4] | proc_20_input_sync_blk[4] | proc_20_output_sync_blk[4]);
    assign proc_20_data_FIFO_blk[5] = 1'b0;
    assign proc_20_data_PIPO_blk[5] = 1'b0;
    assign proc_20_start_FIFO_blk[5] = 1'b0;
    assign proc_20_TLF_FIFO_blk[5] = 1'b0;
    assign proc_20_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_20_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_20[5] = dl_detect_out ? proc_dep_vld_vec_20_reg[5] : (proc_20_data_FIFO_blk[5] | proc_20_data_PIPO_blk[5] | proc_20_start_FIFO_blk[5] | proc_20_TLF_FIFO_blk[5] | proc_20_input_sync_blk[5] | proc_20_output_sync_blk[5]);
    assign proc_20_data_FIFO_blk[6] = 1'b0;
    assign proc_20_data_PIPO_blk[6] = 1'b0;
    assign proc_20_start_FIFO_blk[6] = 1'b0;
    assign proc_20_TLF_FIFO_blk[6] = 1'b0;
    assign proc_20_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_20_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_20[6] = dl_detect_out ? proc_dep_vld_vec_20_reg[6] : (proc_20_data_FIFO_blk[6] | proc_20_data_PIPO_blk[6] | proc_20_start_FIFO_blk[6] | proc_20_TLF_FIFO_blk[6] | proc_20_input_sync_blk[6] | proc_20_output_sync_blk[6]);
    assign proc_20_data_FIFO_blk[7] = 1'b0;
    assign proc_20_data_PIPO_blk[7] = 1'b0;
    assign proc_20_start_FIFO_blk[7] = 1'b0;
    assign proc_20_TLF_FIFO_blk[7] = 1'b0;
    assign proc_20_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_20_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_20[7] = dl_detect_out ? proc_dep_vld_vec_20_reg[7] : (proc_20_data_FIFO_blk[7] | proc_20_data_PIPO_blk[7] | proc_20_start_FIFO_blk[7] | proc_20_TLF_FIFO_blk[7] | proc_20_input_sync_blk[7] | proc_20_output_sync_blk[7]);
    assign proc_20_data_FIFO_blk[8] = 1'b0;
    assign proc_20_data_PIPO_blk[8] = 1'b0;
    assign proc_20_start_FIFO_blk[8] = 1'b0;
    assign proc_20_TLF_FIFO_blk[8] = 1'b0;
    assign proc_20_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_20_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_20[8] = dl_detect_out ? proc_dep_vld_vec_20_reg[8] : (proc_20_data_FIFO_blk[8] | proc_20_data_PIPO_blk[8] | proc_20_start_FIFO_blk[8] | proc_20_TLF_FIFO_blk[8] | proc_20_input_sync_blk[8] | proc_20_output_sync_blk[8]);
    assign proc_20_data_FIFO_blk[9] = 1'b0;
    assign proc_20_data_PIPO_blk[9] = 1'b0;
    assign proc_20_start_FIFO_blk[9] = 1'b0;
    assign proc_20_TLF_FIFO_blk[9] = 1'b0;
    assign proc_20_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_20_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_20[9] = dl_detect_out ? proc_dep_vld_vec_20_reg[9] : (proc_20_data_FIFO_blk[9] | proc_20_data_PIPO_blk[9] | proc_20_start_FIFO_blk[9] | proc_20_TLF_FIFO_blk[9] | proc_20_input_sync_blk[9] | proc_20_output_sync_blk[9]);
    assign proc_20_data_FIFO_blk[10] = 1'b0;
    assign proc_20_data_PIPO_blk[10] = 1'b0;
    assign proc_20_start_FIFO_blk[10] = 1'b0;
    assign proc_20_TLF_FIFO_blk[10] = 1'b0;
    assign proc_20_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_20_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_20[10] = dl_detect_out ? proc_dep_vld_vec_20_reg[10] : (proc_20_data_FIFO_blk[10] | proc_20_data_PIPO_blk[10] | proc_20_start_FIFO_blk[10] | proc_20_TLF_FIFO_blk[10] | proc_20_input_sync_blk[10] | proc_20_output_sync_blk[10]);
    assign proc_20_data_FIFO_blk[11] = 1'b0;
    assign proc_20_data_PIPO_blk[11] = 1'b0;
    assign proc_20_start_FIFO_blk[11] = 1'b0;
    assign proc_20_TLF_FIFO_blk[11] = 1'b0;
    assign proc_20_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_20_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_20[11] = dl_detect_out ? proc_dep_vld_vec_20_reg[11] : (proc_20_data_FIFO_blk[11] | proc_20_data_PIPO_blk[11] | proc_20_start_FIFO_blk[11] | proc_20_TLF_FIFO_blk[11] | proc_20_input_sync_blk[11] | proc_20_output_sync_blk[11]);
    assign proc_20_data_FIFO_blk[12] = 1'b0;
    assign proc_20_data_PIPO_blk[12] = 1'b0;
    assign proc_20_start_FIFO_blk[12] = 1'b0;
    assign proc_20_TLF_FIFO_blk[12] = 1'b0;
    assign proc_20_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_20_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_20[12] = dl_detect_out ? proc_dep_vld_vec_20_reg[12] : (proc_20_data_FIFO_blk[12] | proc_20_data_PIPO_blk[12] | proc_20_start_FIFO_blk[12] | proc_20_TLF_FIFO_blk[12] | proc_20_input_sync_blk[12] | proc_20_output_sync_blk[12]);
    assign proc_20_data_FIFO_blk[13] = 1'b0;
    assign proc_20_data_PIPO_blk[13] = 1'b0;
    assign proc_20_start_FIFO_blk[13] = 1'b0;
    assign proc_20_TLF_FIFO_blk[13] = 1'b0;
    assign proc_20_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_20_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_20[13] = dl_detect_out ? proc_dep_vld_vec_20_reg[13] : (proc_20_data_FIFO_blk[13] | proc_20_data_PIPO_blk[13] | proc_20_start_FIFO_blk[13] | proc_20_TLF_FIFO_blk[13] | proc_20_input_sync_blk[13] | proc_20_output_sync_blk[13]);
    assign proc_20_data_FIFO_blk[14] = 1'b0;
    assign proc_20_data_PIPO_blk[14] = 1'b0;
    assign proc_20_start_FIFO_blk[14] = 1'b0;
    assign proc_20_TLF_FIFO_blk[14] = 1'b0;
    assign proc_20_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_20_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_20[14] = dl_detect_out ? proc_dep_vld_vec_20_reg[14] : (proc_20_data_FIFO_blk[14] | proc_20_data_PIPO_blk[14] | proc_20_start_FIFO_blk[14] | proc_20_TLF_FIFO_blk[14] | proc_20_input_sync_blk[14] | proc_20_output_sync_blk[14]);
    assign proc_20_data_FIFO_blk[15] = 1'b0;
    assign proc_20_data_PIPO_blk[15] = 1'b0;
    assign proc_20_start_FIFO_blk[15] = 1'b0;
    assign proc_20_TLF_FIFO_blk[15] = 1'b0;
    assign proc_20_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_20_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_20[15] = dl_detect_out ? proc_dep_vld_vec_20_reg[15] : (proc_20_data_FIFO_blk[15] | proc_20_data_PIPO_blk[15] | proc_20_start_FIFO_blk[15] | proc_20_TLF_FIFO_blk[15] | proc_20_input_sync_blk[15] | proc_20_output_sync_blk[15]);
    assign proc_20_data_FIFO_blk[16] = 1'b0;
    assign proc_20_data_PIPO_blk[16] = 1'b0;
    assign proc_20_start_FIFO_blk[16] = 1'b0;
    assign proc_20_TLF_FIFO_blk[16] = 1'b0;
    assign proc_20_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_20_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_20[16] = dl_detect_out ? proc_dep_vld_vec_20_reg[16] : (proc_20_data_FIFO_blk[16] | proc_20_data_PIPO_blk[16] | proc_20_start_FIFO_blk[16] | proc_20_TLF_FIFO_blk[16] | proc_20_input_sync_blk[16] | proc_20_output_sync_blk[16]);
    assign proc_20_data_FIFO_blk[17] = 1'b0;
    assign proc_20_data_PIPO_blk[17] = 1'b0;
    assign proc_20_start_FIFO_blk[17] = 1'b0;
    assign proc_20_TLF_FIFO_blk[17] = 1'b0;
    assign proc_20_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_20_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_20[17] = dl_detect_out ? proc_dep_vld_vec_20_reg[17] : (proc_20_data_FIFO_blk[17] | proc_20_data_PIPO_blk[17] | proc_20_start_FIFO_blk[17] | proc_20_TLF_FIFO_blk[17] | proc_20_input_sync_blk[17] | proc_20_output_sync_blk[17]);
    assign proc_20_data_FIFO_blk[18] = 1'b0;
    assign proc_20_data_PIPO_blk[18] = 1'b0;
    assign proc_20_start_FIFO_blk[18] = 1'b0;
    assign proc_20_TLF_FIFO_blk[18] = 1'b0;
    assign proc_20_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_20_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_20[18] = dl_detect_out ? proc_dep_vld_vec_20_reg[18] : (proc_20_data_FIFO_blk[18] | proc_20_data_PIPO_blk[18] | proc_20_start_FIFO_blk[18] | proc_20_TLF_FIFO_blk[18] | proc_20_input_sync_blk[18] | proc_20_output_sync_blk[18]);
    assign proc_20_data_FIFO_blk[19] = 1'b0;
    assign proc_20_data_PIPO_blk[19] = 1'b0;
    assign proc_20_start_FIFO_blk[19] = 1'b0;
    assign proc_20_TLF_FIFO_blk[19] = 1'b0;
    assign proc_20_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_20_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_20[19] = dl_detect_out ? proc_dep_vld_vec_20_reg[19] : (proc_20_data_FIFO_blk[19] | proc_20_data_PIPO_blk[19] | proc_20_start_FIFO_blk[19] | proc_20_TLF_FIFO_blk[19] | proc_20_input_sync_blk[19] | proc_20_output_sync_blk[19]);
    assign proc_20_data_FIFO_blk[20] = 1'b0;
    assign proc_20_data_PIPO_blk[20] = 1'b0;
    assign proc_20_start_FIFO_blk[20] = 1'b0;
    assign proc_20_TLF_FIFO_blk[20] = 1'b0;
    assign proc_20_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_20_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_20[20] = dl_detect_out ? proc_dep_vld_vec_20_reg[20] : (proc_20_data_FIFO_blk[20] | proc_20_data_PIPO_blk[20] | proc_20_start_FIFO_blk[20] | proc_20_TLF_FIFO_blk[20] | proc_20_input_sync_blk[20] | proc_20_output_sync_blk[20]);
    assign proc_20_data_FIFO_blk[21] = 1'b0;
    assign proc_20_data_PIPO_blk[21] = 1'b0;
    assign proc_20_start_FIFO_blk[21] = 1'b0;
    assign proc_20_TLF_FIFO_blk[21] = 1'b0;
    assign proc_20_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_20_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_20[21] = dl_detect_out ? proc_dep_vld_vec_20_reg[21] : (proc_20_data_FIFO_blk[21] | proc_20_data_PIPO_blk[21] | proc_20_start_FIFO_blk[21] | proc_20_TLF_FIFO_blk[21] | proc_20_input_sync_blk[21] | proc_20_output_sync_blk[21]);
    assign proc_20_data_FIFO_blk[22] = 1'b0;
    assign proc_20_data_PIPO_blk[22] = 1'b0;
    assign proc_20_start_FIFO_blk[22] = 1'b0;
    assign proc_20_TLF_FIFO_blk[22] = 1'b0;
    assign proc_20_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_20_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_20[22] = dl_detect_out ? proc_dep_vld_vec_20_reg[22] : (proc_20_data_FIFO_blk[22] | proc_20_data_PIPO_blk[22] | proc_20_start_FIFO_blk[22] | proc_20_TLF_FIFO_blk[22] | proc_20_input_sync_blk[22] | proc_20_output_sync_blk[22]);
    assign proc_20_data_FIFO_blk[23] = 1'b0;
    assign proc_20_data_PIPO_blk[23] = 1'b0;
    assign proc_20_start_FIFO_blk[23] = 1'b0;
    assign proc_20_TLF_FIFO_blk[23] = 1'b0;
    assign proc_20_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_20_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_20[23] = dl_detect_out ? proc_dep_vld_vec_20_reg[23] : (proc_20_data_FIFO_blk[23] | proc_20_data_PIPO_blk[23] | proc_20_start_FIFO_blk[23] | proc_20_TLF_FIFO_blk[23] | proc_20_input_sync_blk[23] | proc_20_output_sync_blk[23]);
    assign proc_20_data_FIFO_blk[24] = 1'b0;
    assign proc_20_data_PIPO_blk[24] = 1'b0;
    assign proc_20_start_FIFO_blk[24] = 1'b0;
    assign proc_20_TLF_FIFO_blk[24] = 1'b0;
    assign proc_20_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_20_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_20[24] = dl_detect_out ? proc_dep_vld_vec_20_reg[24] : (proc_20_data_FIFO_blk[24] | proc_20_data_PIPO_blk[24] | proc_20_start_FIFO_blk[24] | proc_20_TLF_FIFO_blk[24] | proc_20_input_sync_blk[24] | proc_20_output_sync_blk[24]);
    assign proc_20_data_FIFO_blk[25] = 1'b0;
    assign proc_20_data_PIPO_blk[25] = 1'b0;
    assign proc_20_start_FIFO_blk[25] = 1'b0;
    assign proc_20_TLF_FIFO_blk[25] = 1'b0;
    assign proc_20_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_20_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_20[25] = dl_detect_out ? proc_dep_vld_vec_20_reg[25] : (proc_20_data_FIFO_blk[25] | proc_20_data_PIPO_blk[25] | proc_20_start_FIFO_blk[25] | proc_20_TLF_FIFO_blk[25] | proc_20_input_sync_blk[25] | proc_20_output_sync_blk[25]);
    assign proc_20_data_FIFO_blk[26] = 1'b0;
    assign proc_20_data_PIPO_blk[26] = 1'b0;
    assign proc_20_start_FIFO_blk[26] = 1'b0;
    assign proc_20_TLF_FIFO_blk[26] = 1'b0;
    assign proc_20_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_20_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_20[26] = dl_detect_out ? proc_dep_vld_vec_20_reg[26] : (proc_20_data_FIFO_blk[26] | proc_20_data_PIPO_blk[26] | proc_20_start_FIFO_blk[26] | proc_20_TLF_FIFO_blk[26] | proc_20_input_sync_blk[26] | proc_20_output_sync_blk[26]);
    assign proc_20_data_FIFO_blk[27] = 1'b0;
    assign proc_20_data_PIPO_blk[27] = 1'b0;
    assign proc_20_start_FIFO_blk[27] = 1'b0;
    assign proc_20_TLF_FIFO_blk[27] = 1'b0;
    assign proc_20_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_20_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_20[27] = dl_detect_out ? proc_dep_vld_vec_20_reg[27] : (proc_20_data_FIFO_blk[27] | proc_20_data_PIPO_blk[27] | proc_20_start_FIFO_blk[27] | proc_20_TLF_FIFO_blk[27] | proc_20_input_sync_blk[27] | proc_20_output_sync_blk[27]);
    assign proc_20_data_FIFO_blk[28] = 1'b0;
    assign proc_20_data_PIPO_blk[28] = 1'b0;
    assign proc_20_start_FIFO_blk[28] = 1'b0;
    assign proc_20_TLF_FIFO_blk[28] = 1'b0;
    assign proc_20_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_20_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_20[28] = dl_detect_out ? proc_dep_vld_vec_20_reg[28] : (proc_20_data_FIFO_blk[28] | proc_20_data_PIPO_blk[28] | proc_20_start_FIFO_blk[28] | proc_20_TLF_FIFO_blk[28] | proc_20_input_sync_blk[28] | proc_20_output_sync_blk[28]);
    assign proc_20_data_FIFO_blk[29] = 1'b0;
    assign proc_20_data_PIPO_blk[29] = 1'b0;
    assign proc_20_start_FIFO_blk[29] = 1'b0;
    assign proc_20_TLF_FIFO_blk[29] = 1'b0;
    assign proc_20_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_20_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_20[29] = dl_detect_out ? proc_dep_vld_vec_20_reg[29] : (proc_20_data_FIFO_blk[29] | proc_20_data_PIPO_blk[29] | proc_20_start_FIFO_blk[29] | proc_20_TLF_FIFO_blk[29] | proc_20_input_sync_blk[29] | proc_20_output_sync_blk[29]);
    assign proc_20_data_FIFO_blk[30] = 1'b0;
    assign proc_20_data_PIPO_blk[30] = 1'b0;
    assign proc_20_start_FIFO_blk[30] = 1'b0;
    assign proc_20_TLF_FIFO_blk[30] = 1'b0;
    assign proc_20_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_20_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_20[30] = dl_detect_out ? proc_dep_vld_vec_20_reg[30] : (proc_20_data_FIFO_blk[30] | proc_20_data_PIPO_blk[30] | proc_20_start_FIFO_blk[30] | proc_20_TLF_FIFO_blk[30] | proc_20_input_sync_blk[30] | proc_20_output_sync_blk[30]);
    assign proc_20_data_FIFO_blk[31] = 1'b0;
    assign proc_20_data_PIPO_blk[31] = 1'b0;
    assign proc_20_start_FIFO_blk[31] = 1'b0;
    assign proc_20_TLF_FIFO_blk[31] = 1'b0;
    assign proc_20_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_20_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_20[31] = dl_detect_out ? proc_dep_vld_vec_20_reg[31] : (proc_20_data_FIFO_blk[31] | proc_20_data_PIPO_blk[31] | proc_20_start_FIFO_blk[31] | proc_20_TLF_FIFO_blk[31] | proc_20_input_sync_blk[31] | proc_20_output_sync_blk[31]);
    assign proc_20_data_FIFO_blk[32] = 1'b0;
    assign proc_20_data_PIPO_blk[32] = 1'b0;
    assign proc_20_start_FIFO_blk[32] = 1'b0;
    assign proc_20_TLF_FIFO_blk[32] = 1'b0;
    assign proc_20_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_15_U0_ap_ready & ProcessingElement_15_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_20_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_20[32] = dl_detect_out ? proc_dep_vld_vec_20_reg[32] : (proc_20_data_FIFO_blk[32] | proc_20_data_PIPO_blk[32] | proc_20_start_FIFO_blk[32] | proc_20_TLF_FIFO_blk[32] | proc_20_input_sync_blk[32] | proc_20_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_20_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_20_reg <= proc_dep_vld_vec_20;
        end
    end
    assign in_chan_dep_vld_vec_20[0] = dep_chan_vld_0_20;
    assign in_chan_dep_data_vec_20[39 : 0] = dep_chan_data_0_20;
    assign token_in_vec_20[0] = token_0_20;
    assign in_chan_dep_vld_vec_20[1] = dep_chan_vld_1_20;
    assign in_chan_dep_data_vec_20[79 : 40] = dep_chan_data_1_20;
    assign token_in_vec_20[1] = token_1_20;
    assign in_chan_dep_vld_vec_20[2] = dep_chan_vld_3_20;
    assign in_chan_dep_data_vec_20[119 : 80] = dep_chan_data_3_20;
    assign token_in_vec_20[2] = token_3_20;
    assign in_chan_dep_vld_vec_20[3] = dep_chan_vld_6_20;
    assign in_chan_dep_data_vec_20[159 : 120] = dep_chan_data_6_20;
    assign token_in_vec_20[3] = token_6_20;
    assign in_chan_dep_vld_vec_20[4] = dep_chan_vld_7_20;
    assign in_chan_dep_data_vec_20[199 : 160] = dep_chan_data_7_20;
    assign token_in_vec_20[4] = token_7_20;
    assign in_chan_dep_vld_vec_20[5] = dep_chan_vld_8_20;
    assign in_chan_dep_data_vec_20[239 : 200] = dep_chan_data_8_20;
    assign token_in_vec_20[5] = token_8_20;
    assign in_chan_dep_vld_vec_20[6] = dep_chan_vld_9_20;
    assign in_chan_dep_data_vec_20[279 : 240] = dep_chan_data_9_20;
    assign token_in_vec_20[6] = token_9_20;
    assign in_chan_dep_vld_vec_20[7] = dep_chan_vld_10_20;
    assign in_chan_dep_data_vec_20[319 : 280] = dep_chan_data_10_20;
    assign token_in_vec_20[7] = token_10_20;
    assign in_chan_dep_vld_vec_20[8] = dep_chan_vld_11_20;
    assign in_chan_dep_data_vec_20[359 : 320] = dep_chan_data_11_20;
    assign token_in_vec_20[8] = token_11_20;
    assign in_chan_dep_vld_vec_20[9] = dep_chan_vld_12_20;
    assign in_chan_dep_data_vec_20[399 : 360] = dep_chan_data_12_20;
    assign token_in_vec_20[9] = token_12_20;
    assign in_chan_dep_vld_vec_20[10] = dep_chan_vld_13_20;
    assign in_chan_dep_data_vec_20[439 : 400] = dep_chan_data_13_20;
    assign token_in_vec_20[10] = token_13_20;
    assign in_chan_dep_vld_vec_20[11] = dep_chan_vld_14_20;
    assign in_chan_dep_data_vec_20[479 : 440] = dep_chan_data_14_20;
    assign token_in_vec_20[11] = token_14_20;
    assign in_chan_dep_vld_vec_20[12] = dep_chan_vld_15_20;
    assign in_chan_dep_data_vec_20[519 : 480] = dep_chan_data_15_20;
    assign token_in_vec_20[12] = token_15_20;
    assign in_chan_dep_vld_vec_20[13] = dep_chan_vld_16_20;
    assign in_chan_dep_data_vec_20[559 : 520] = dep_chan_data_16_20;
    assign token_in_vec_20[13] = token_16_20;
    assign in_chan_dep_vld_vec_20[14] = dep_chan_vld_17_20;
    assign in_chan_dep_data_vec_20[599 : 560] = dep_chan_data_17_20;
    assign token_in_vec_20[14] = token_17_20;
    assign in_chan_dep_vld_vec_20[15] = dep_chan_vld_18_20;
    assign in_chan_dep_data_vec_20[639 : 600] = dep_chan_data_18_20;
    assign token_in_vec_20[15] = token_18_20;
    assign in_chan_dep_vld_vec_20[16] = dep_chan_vld_19_20;
    assign in_chan_dep_data_vec_20[679 : 640] = dep_chan_data_19_20;
    assign token_in_vec_20[16] = token_19_20;
    assign in_chan_dep_vld_vec_20[17] = dep_chan_vld_21_20;
    assign in_chan_dep_data_vec_20[719 : 680] = dep_chan_data_21_20;
    assign token_in_vec_20[17] = token_21_20;
    assign in_chan_dep_vld_vec_20[18] = dep_chan_vld_22_20;
    assign in_chan_dep_data_vec_20[759 : 720] = dep_chan_data_22_20;
    assign token_in_vec_20[18] = token_22_20;
    assign in_chan_dep_vld_vec_20[19] = dep_chan_vld_23_20;
    assign in_chan_dep_data_vec_20[799 : 760] = dep_chan_data_23_20;
    assign token_in_vec_20[19] = token_23_20;
    assign in_chan_dep_vld_vec_20[20] = dep_chan_vld_24_20;
    assign in_chan_dep_data_vec_20[839 : 800] = dep_chan_data_24_20;
    assign token_in_vec_20[20] = token_24_20;
    assign in_chan_dep_vld_vec_20[21] = dep_chan_vld_25_20;
    assign in_chan_dep_data_vec_20[879 : 840] = dep_chan_data_25_20;
    assign token_in_vec_20[21] = token_25_20;
    assign in_chan_dep_vld_vec_20[22] = dep_chan_vld_26_20;
    assign in_chan_dep_data_vec_20[919 : 880] = dep_chan_data_26_20;
    assign token_in_vec_20[22] = token_26_20;
    assign in_chan_dep_vld_vec_20[23] = dep_chan_vld_27_20;
    assign in_chan_dep_data_vec_20[959 : 920] = dep_chan_data_27_20;
    assign token_in_vec_20[23] = token_27_20;
    assign in_chan_dep_vld_vec_20[24] = dep_chan_vld_28_20;
    assign in_chan_dep_data_vec_20[999 : 960] = dep_chan_data_28_20;
    assign token_in_vec_20[24] = token_28_20;
    assign in_chan_dep_vld_vec_20[25] = dep_chan_vld_29_20;
    assign in_chan_dep_data_vec_20[1039 : 1000] = dep_chan_data_29_20;
    assign token_in_vec_20[25] = token_29_20;
    assign in_chan_dep_vld_vec_20[26] = dep_chan_vld_30_20;
    assign in_chan_dep_data_vec_20[1079 : 1040] = dep_chan_data_30_20;
    assign token_in_vec_20[26] = token_30_20;
    assign in_chan_dep_vld_vec_20[27] = dep_chan_vld_31_20;
    assign in_chan_dep_data_vec_20[1119 : 1080] = dep_chan_data_31_20;
    assign token_in_vec_20[27] = token_31_20;
    assign in_chan_dep_vld_vec_20[28] = dep_chan_vld_32_20;
    assign in_chan_dep_data_vec_20[1159 : 1120] = dep_chan_data_32_20;
    assign token_in_vec_20[28] = token_32_20;
    assign in_chan_dep_vld_vec_20[29] = dep_chan_vld_33_20;
    assign in_chan_dep_data_vec_20[1199 : 1160] = dep_chan_data_33_20;
    assign token_in_vec_20[29] = token_33_20;
    assign in_chan_dep_vld_vec_20[30] = dep_chan_vld_34_20;
    assign in_chan_dep_data_vec_20[1239 : 1200] = dep_chan_data_34_20;
    assign token_in_vec_20[30] = token_34_20;
    assign in_chan_dep_vld_vec_20[31] = dep_chan_vld_35_20;
    assign in_chan_dep_data_vec_20[1279 : 1240] = dep_chan_data_35_20;
    assign token_in_vec_20[31] = token_35_20;
    assign in_chan_dep_vld_vec_20[32] = dep_chan_vld_36_20;
    assign in_chan_dep_data_vec_20[1319 : 1280] = dep_chan_data_36_20;
    assign token_in_vec_20[32] = token_36_20;
    assign dep_chan_vld_20_19 = out_chan_dep_vld_vec_20[0];
    assign dep_chan_data_20_19 = out_chan_dep_data_20;
    assign token_20_19 = token_out_vec_20[0];
    assign dep_chan_vld_20_21 = out_chan_dep_vld_vec_20[1];
    assign dep_chan_data_20_21 = out_chan_dep_data_20;
    assign token_20_21 = token_out_vec_20[1];
    assign dep_chan_vld_20_0 = out_chan_dep_vld_vec_20[2];
    assign dep_chan_data_20_0 = out_chan_dep_data_20;
    assign token_20_0 = token_out_vec_20[2];
    assign dep_chan_vld_20_1 = out_chan_dep_vld_vec_20[3];
    assign dep_chan_data_20_1 = out_chan_dep_data_20;
    assign token_20_1 = token_out_vec_20[3];
    assign dep_chan_vld_20_3 = out_chan_dep_vld_vec_20[4];
    assign dep_chan_data_20_3 = out_chan_dep_data_20;
    assign token_20_3 = token_out_vec_20[4];
    assign dep_chan_vld_20_6 = out_chan_dep_vld_vec_20[5];
    assign dep_chan_data_20_6 = out_chan_dep_data_20;
    assign token_20_6 = token_out_vec_20[5];
    assign dep_chan_vld_20_7 = out_chan_dep_vld_vec_20[6];
    assign dep_chan_data_20_7 = out_chan_dep_data_20;
    assign token_20_7 = token_out_vec_20[6];
    assign dep_chan_vld_20_8 = out_chan_dep_vld_vec_20[7];
    assign dep_chan_data_20_8 = out_chan_dep_data_20;
    assign token_20_8 = token_out_vec_20[7];
    assign dep_chan_vld_20_9 = out_chan_dep_vld_vec_20[8];
    assign dep_chan_data_20_9 = out_chan_dep_data_20;
    assign token_20_9 = token_out_vec_20[8];
    assign dep_chan_vld_20_10 = out_chan_dep_vld_vec_20[9];
    assign dep_chan_data_20_10 = out_chan_dep_data_20;
    assign token_20_10 = token_out_vec_20[9];
    assign dep_chan_vld_20_11 = out_chan_dep_vld_vec_20[10];
    assign dep_chan_data_20_11 = out_chan_dep_data_20;
    assign token_20_11 = token_out_vec_20[10];
    assign dep_chan_vld_20_12 = out_chan_dep_vld_vec_20[11];
    assign dep_chan_data_20_12 = out_chan_dep_data_20;
    assign token_20_12 = token_out_vec_20[11];
    assign dep_chan_vld_20_13 = out_chan_dep_vld_vec_20[12];
    assign dep_chan_data_20_13 = out_chan_dep_data_20;
    assign token_20_13 = token_out_vec_20[12];
    assign dep_chan_vld_20_14 = out_chan_dep_vld_vec_20[13];
    assign dep_chan_data_20_14 = out_chan_dep_data_20;
    assign token_20_14 = token_out_vec_20[13];
    assign dep_chan_vld_20_15 = out_chan_dep_vld_vec_20[14];
    assign dep_chan_data_20_15 = out_chan_dep_data_20;
    assign token_20_15 = token_out_vec_20[14];
    assign dep_chan_vld_20_16 = out_chan_dep_vld_vec_20[15];
    assign dep_chan_data_20_16 = out_chan_dep_data_20;
    assign token_20_16 = token_out_vec_20[15];
    assign dep_chan_vld_20_17 = out_chan_dep_vld_vec_20[16];
    assign dep_chan_data_20_17 = out_chan_dep_data_20;
    assign token_20_17 = token_out_vec_20[16];
    assign dep_chan_vld_20_18 = out_chan_dep_vld_vec_20[17];
    assign dep_chan_data_20_18 = out_chan_dep_data_20;
    assign token_20_18 = token_out_vec_20[17];
    assign dep_chan_vld_20_22 = out_chan_dep_vld_vec_20[18];
    assign dep_chan_data_20_22 = out_chan_dep_data_20;
    assign token_20_22 = token_out_vec_20[18];
    assign dep_chan_vld_20_23 = out_chan_dep_vld_vec_20[19];
    assign dep_chan_data_20_23 = out_chan_dep_data_20;
    assign token_20_23 = token_out_vec_20[19];
    assign dep_chan_vld_20_24 = out_chan_dep_vld_vec_20[20];
    assign dep_chan_data_20_24 = out_chan_dep_data_20;
    assign token_20_24 = token_out_vec_20[20];
    assign dep_chan_vld_20_25 = out_chan_dep_vld_vec_20[21];
    assign dep_chan_data_20_25 = out_chan_dep_data_20;
    assign token_20_25 = token_out_vec_20[21];
    assign dep_chan_vld_20_26 = out_chan_dep_vld_vec_20[22];
    assign dep_chan_data_20_26 = out_chan_dep_data_20;
    assign token_20_26 = token_out_vec_20[22];
    assign dep_chan_vld_20_27 = out_chan_dep_vld_vec_20[23];
    assign dep_chan_data_20_27 = out_chan_dep_data_20;
    assign token_20_27 = token_out_vec_20[23];
    assign dep_chan_vld_20_28 = out_chan_dep_vld_vec_20[24];
    assign dep_chan_data_20_28 = out_chan_dep_data_20;
    assign token_20_28 = token_out_vec_20[24];
    assign dep_chan_vld_20_29 = out_chan_dep_vld_vec_20[25];
    assign dep_chan_data_20_29 = out_chan_dep_data_20;
    assign token_20_29 = token_out_vec_20[25];
    assign dep_chan_vld_20_30 = out_chan_dep_vld_vec_20[26];
    assign dep_chan_data_20_30 = out_chan_dep_data_20;
    assign token_20_30 = token_out_vec_20[26];
    assign dep_chan_vld_20_31 = out_chan_dep_vld_vec_20[27];
    assign dep_chan_data_20_31 = out_chan_dep_data_20;
    assign token_20_31 = token_out_vec_20[27];
    assign dep_chan_vld_20_32 = out_chan_dep_vld_vec_20[28];
    assign dep_chan_data_20_32 = out_chan_dep_data_20;
    assign token_20_32 = token_out_vec_20[28];
    assign dep_chan_vld_20_33 = out_chan_dep_vld_vec_20[29];
    assign dep_chan_data_20_33 = out_chan_dep_data_20;
    assign token_20_33 = token_out_vec_20[29];
    assign dep_chan_vld_20_34 = out_chan_dep_vld_vec_20[30];
    assign dep_chan_data_20_34 = out_chan_dep_data_20;
    assign token_20_34 = token_out_vec_20[30];
    assign dep_chan_vld_20_35 = out_chan_dep_vld_vec_20[31];
    assign dep_chan_data_20_35 = out_chan_dep_data_20;
    assign token_20_35 = token_out_vec_20[31];
    assign dep_chan_vld_20_36 = out_chan_dep_vld_vec_20[32];
    assign dep_chan_data_20_36 = out_chan_dep_data_20;
    assign token_20_36 = token_out_vec_20[32];

    // Process: ProcessingElement_16_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 21, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_21 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_21),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_21),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_21),
        .token_in_vec(token_in_vec_21),
        .dl_detect_in(dl_detect_out),
        .origin(origin[21]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_21),
        .out_chan_dep_data(out_chan_dep_data_21),
        .token_out_vec(token_out_vec_21),
        .dl_detect_out(dl_in_vec[21]));

    assign proc_21_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_15_blk_n) | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_15_blk_n) | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_WriteC_Flattened_fu_179.cPipes_15_blk_n);
    assign proc_21_data_PIPO_blk[0] = 1'b0;
    assign proc_21_start_FIFO_blk[0] = 1'b0;
    assign proc_21_TLF_FIFO_blk[0] = 1'b0;
    assign proc_21_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_21_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_21[0] = dl_detect_out ? proc_dep_vld_vec_21_reg[0] : (proc_21_data_FIFO_blk[0] | proc_21_data_PIPO_blk[0] | proc_21_start_FIFO_blk[0] | proc_21_TLF_FIFO_blk[0] | proc_21_input_sync_blk[0] | proc_21_output_sync_blk[0]);
    assign proc_21_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_16_blk_n) | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_16_blk_n) | (~ProcessingElement_16_U0.grp_ProcessingElement_16_Pipeline_WriteC_Flattened_fu_179.cPipes_16_blk_n);
    assign proc_21_data_PIPO_blk[1] = 1'b0;
    assign proc_21_start_FIFO_blk[1] = 1'b0;
    assign proc_21_TLF_FIFO_blk[1] = 1'b0;
    assign proc_21_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_21_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_21[1] = dl_detect_out ? proc_dep_vld_vec_21_reg[1] : (proc_21_data_FIFO_blk[1] | proc_21_data_PIPO_blk[1] | proc_21_start_FIFO_blk[1] | proc_21_TLF_FIFO_blk[1] | proc_21_input_sync_blk[1] | proc_21_output_sync_blk[1]);
    assign proc_21_data_FIFO_blk[2] = 1'b0;
    assign proc_21_data_PIPO_blk[2] = 1'b0;
    assign proc_21_start_FIFO_blk[2] = 1'b0;
    assign proc_21_TLF_FIFO_blk[2] = 1'b0;
    assign proc_21_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_21_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_21[2] = dl_detect_out ? proc_dep_vld_vec_21_reg[2] : (proc_21_data_FIFO_blk[2] | proc_21_data_PIPO_blk[2] | proc_21_start_FIFO_blk[2] | proc_21_TLF_FIFO_blk[2] | proc_21_input_sync_blk[2] | proc_21_output_sync_blk[2]);
    assign proc_21_data_FIFO_blk[3] = 1'b0;
    assign proc_21_data_PIPO_blk[3] = 1'b0;
    assign proc_21_start_FIFO_blk[3] = 1'b0;
    assign proc_21_TLF_FIFO_blk[3] = 1'b0;
    assign proc_21_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_21_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_21[3] = dl_detect_out ? proc_dep_vld_vec_21_reg[3] : (proc_21_data_FIFO_blk[3] | proc_21_data_PIPO_blk[3] | proc_21_start_FIFO_blk[3] | proc_21_TLF_FIFO_blk[3] | proc_21_input_sync_blk[3] | proc_21_output_sync_blk[3]);
    assign proc_21_data_FIFO_blk[4] = 1'b0;
    assign proc_21_data_PIPO_blk[4] = 1'b0;
    assign proc_21_start_FIFO_blk[4] = 1'b0;
    assign proc_21_TLF_FIFO_blk[4] = 1'b0;
    assign proc_21_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_21_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_21[4] = dl_detect_out ? proc_dep_vld_vec_21_reg[4] : (proc_21_data_FIFO_blk[4] | proc_21_data_PIPO_blk[4] | proc_21_start_FIFO_blk[4] | proc_21_TLF_FIFO_blk[4] | proc_21_input_sync_blk[4] | proc_21_output_sync_blk[4]);
    assign proc_21_data_FIFO_blk[5] = 1'b0;
    assign proc_21_data_PIPO_blk[5] = 1'b0;
    assign proc_21_start_FIFO_blk[5] = 1'b0;
    assign proc_21_TLF_FIFO_blk[5] = 1'b0;
    assign proc_21_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_21_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_21[5] = dl_detect_out ? proc_dep_vld_vec_21_reg[5] : (proc_21_data_FIFO_blk[5] | proc_21_data_PIPO_blk[5] | proc_21_start_FIFO_blk[5] | proc_21_TLF_FIFO_blk[5] | proc_21_input_sync_blk[5] | proc_21_output_sync_blk[5]);
    assign proc_21_data_FIFO_blk[6] = 1'b0;
    assign proc_21_data_PIPO_blk[6] = 1'b0;
    assign proc_21_start_FIFO_blk[6] = 1'b0;
    assign proc_21_TLF_FIFO_blk[6] = 1'b0;
    assign proc_21_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_21_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_21[6] = dl_detect_out ? proc_dep_vld_vec_21_reg[6] : (proc_21_data_FIFO_blk[6] | proc_21_data_PIPO_blk[6] | proc_21_start_FIFO_blk[6] | proc_21_TLF_FIFO_blk[6] | proc_21_input_sync_blk[6] | proc_21_output_sync_blk[6]);
    assign proc_21_data_FIFO_blk[7] = 1'b0;
    assign proc_21_data_PIPO_blk[7] = 1'b0;
    assign proc_21_start_FIFO_blk[7] = 1'b0;
    assign proc_21_TLF_FIFO_blk[7] = 1'b0;
    assign proc_21_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_21_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_21[7] = dl_detect_out ? proc_dep_vld_vec_21_reg[7] : (proc_21_data_FIFO_blk[7] | proc_21_data_PIPO_blk[7] | proc_21_start_FIFO_blk[7] | proc_21_TLF_FIFO_blk[7] | proc_21_input_sync_blk[7] | proc_21_output_sync_blk[7]);
    assign proc_21_data_FIFO_blk[8] = 1'b0;
    assign proc_21_data_PIPO_blk[8] = 1'b0;
    assign proc_21_start_FIFO_blk[8] = 1'b0;
    assign proc_21_TLF_FIFO_blk[8] = 1'b0;
    assign proc_21_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_21_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_21[8] = dl_detect_out ? proc_dep_vld_vec_21_reg[8] : (proc_21_data_FIFO_blk[8] | proc_21_data_PIPO_blk[8] | proc_21_start_FIFO_blk[8] | proc_21_TLF_FIFO_blk[8] | proc_21_input_sync_blk[8] | proc_21_output_sync_blk[8]);
    assign proc_21_data_FIFO_blk[9] = 1'b0;
    assign proc_21_data_PIPO_blk[9] = 1'b0;
    assign proc_21_start_FIFO_blk[9] = 1'b0;
    assign proc_21_TLF_FIFO_blk[9] = 1'b0;
    assign proc_21_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_21_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_21[9] = dl_detect_out ? proc_dep_vld_vec_21_reg[9] : (proc_21_data_FIFO_blk[9] | proc_21_data_PIPO_blk[9] | proc_21_start_FIFO_blk[9] | proc_21_TLF_FIFO_blk[9] | proc_21_input_sync_blk[9] | proc_21_output_sync_blk[9]);
    assign proc_21_data_FIFO_blk[10] = 1'b0;
    assign proc_21_data_PIPO_blk[10] = 1'b0;
    assign proc_21_start_FIFO_blk[10] = 1'b0;
    assign proc_21_TLF_FIFO_blk[10] = 1'b0;
    assign proc_21_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_21_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_21[10] = dl_detect_out ? proc_dep_vld_vec_21_reg[10] : (proc_21_data_FIFO_blk[10] | proc_21_data_PIPO_blk[10] | proc_21_start_FIFO_blk[10] | proc_21_TLF_FIFO_blk[10] | proc_21_input_sync_blk[10] | proc_21_output_sync_blk[10]);
    assign proc_21_data_FIFO_blk[11] = 1'b0;
    assign proc_21_data_PIPO_blk[11] = 1'b0;
    assign proc_21_start_FIFO_blk[11] = 1'b0;
    assign proc_21_TLF_FIFO_blk[11] = 1'b0;
    assign proc_21_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_21_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_21[11] = dl_detect_out ? proc_dep_vld_vec_21_reg[11] : (proc_21_data_FIFO_blk[11] | proc_21_data_PIPO_blk[11] | proc_21_start_FIFO_blk[11] | proc_21_TLF_FIFO_blk[11] | proc_21_input_sync_blk[11] | proc_21_output_sync_blk[11]);
    assign proc_21_data_FIFO_blk[12] = 1'b0;
    assign proc_21_data_PIPO_blk[12] = 1'b0;
    assign proc_21_start_FIFO_blk[12] = 1'b0;
    assign proc_21_TLF_FIFO_blk[12] = 1'b0;
    assign proc_21_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_21_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_21[12] = dl_detect_out ? proc_dep_vld_vec_21_reg[12] : (proc_21_data_FIFO_blk[12] | proc_21_data_PIPO_blk[12] | proc_21_start_FIFO_blk[12] | proc_21_TLF_FIFO_blk[12] | proc_21_input_sync_blk[12] | proc_21_output_sync_blk[12]);
    assign proc_21_data_FIFO_blk[13] = 1'b0;
    assign proc_21_data_PIPO_blk[13] = 1'b0;
    assign proc_21_start_FIFO_blk[13] = 1'b0;
    assign proc_21_TLF_FIFO_blk[13] = 1'b0;
    assign proc_21_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_21_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_21[13] = dl_detect_out ? proc_dep_vld_vec_21_reg[13] : (proc_21_data_FIFO_blk[13] | proc_21_data_PIPO_blk[13] | proc_21_start_FIFO_blk[13] | proc_21_TLF_FIFO_blk[13] | proc_21_input_sync_blk[13] | proc_21_output_sync_blk[13]);
    assign proc_21_data_FIFO_blk[14] = 1'b0;
    assign proc_21_data_PIPO_blk[14] = 1'b0;
    assign proc_21_start_FIFO_blk[14] = 1'b0;
    assign proc_21_TLF_FIFO_blk[14] = 1'b0;
    assign proc_21_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_21_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_21[14] = dl_detect_out ? proc_dep_vld_vec_21_reg[14] : (proc_21_data_FIFO_blk[14] | proc_21_data_PIPO_blk[14] | proc_21_start_FIFO_blk[14] | proc_21_TLF_FIFO_blk[14] | proc_21_input_sync_blk[14] | proc_21_output_sync_blk[14]);
    assign proc_21_data_FIFO_blk[15] = 1'b0;
    assign proc_21_data_PIPO_blk[15] = 1'b0;
    assign proc_21_start_FIFO_blk[15] = 1'b0;
    assign proc_21_TLF_FIFO_blk[15] = 1'b0;
    assign proc_21_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_21_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_21[15] = dl_detect_out ? proc_dep_vld_vec_21_reg[15] : (proc_21_data_FIFO_blk[15] | proc_21_data_PIPO_blk[15] | proc_21_start_FIFO_blk[15] | proc_21_TLF_FIFO_blk[15] | proc_21_input_sync_blk[15] | proc_21_output_sync_blk[15]);
    assign proc_21_data_FIFO_blk[16] = 1'b0;
    assign proc_21_data_PIPO_blk[16] = 1'b0;
    assign proc_21_start_FIFO_blk[16] = 1'b0;
    assign proc_21_TLF_FIFO_blk[16] = 1'b0;
    assign proc_21_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_21_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_21[16] = dl_detect_out ? proc_dep_vld_vec_21_reg[16] : (proc_21_data_FIFO_blk[16] | proc_21_data_PIPO_blk[16] | proc_21_start_FIFO_blk[16] | proc_21_TLF_FIFO_blk[16] | proc_21_input_sync_blk[16] | proc_21_output_sync_blk[16]);
    assign proc_21_data_FIFO_blk[17] = 1'b0;
    assign proc_21_data_PIPO_blk[17] = 1'b0;
    assign proc_21_start_FIFO_blk[17] = 1'b0;
    assign proc_21_TLF_FIFO_blk[17] = 1'b0;
    assign proc_21_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_21_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_21[17] = dl_detect_out ? proc_dep_vld_vec_21_reg[17] : (proc_21_data_FIFO_blk[17] | proc_21_data_PIPO_blk[17] | proc_21_start_FIFO_blk[17] | proc_21_TLF_FIFO_blk[17] | proc_21_input_sync_blk[17] | proc_21_output_sync_blk[17]);
    assign proc_21_data_FIFO_blk[18] = 1'b0;
    assign proc_21_data_PIPO_blk[18] = 1'b0;
    assign proc_21_start_FIFO_blk[18] = 1'b0;
    assign proc_21_TLF_FIFO_blk[18] = 1'b0;
    assign proc_21_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_21_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_21[18] = dl_detect_out ? proc_dep_vld_vec_21_reg[18] : (proc_21_data_FIFO_blk[18] | proc_21_data_PIPO_blk[18] | proc_21_start_FIFO_blk[18] | proc_21_TLF_FIFO_blk[18] | proc_21_input_sync_blk[18] | proc_21_output_sync_blk[18]);
    assign proc_21_data_FIFO_blk[19] = 1'b0;
    assign proc_21_data_PIPO_blk[19] = 1'b0;
    assign proc_21_start_FIFO_blk[19] = 1'b0;
    assign proc_21_TLF_FIFO_blk[19] = 1'b0;
    assign proc_21_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_21_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_21[19] = dl_detect_out ? proc_dep_vld_vec_21_reg[19] : (proc_21_data_FIFO_blk[19] | proc_21_data_PIPO_blk[19] | proc_21_start_FIFO_blk[19] | proc_21_TLF_FIFO_blk[19] | proc_21_input_sync_blk[19] | proc_21_output_sync_blk[19]);
    assign proc_21_data_FIFO_blk[20] = 1'b0;
    assign proc_21_data_PIPO_blk[20] = 1'b0;
    assign proc_21_start_FIFO_blk[20] = 1'b0;
    assign proc_21_TLF_FIFO_blk[20] = 1'b0;
    assign proc_21_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_21_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_21[20] = dl_detect_out ? proc_dep_vld_vec_21_reg[20] : (proc_21_data_FIFO_blk[20] | proc_21_data_PIPO_blk[20] | proc_21_start_FIFO_blk[20] | proc_21_TLF_FIFO_blk[20] | proc_21_input_sync_blk[20] | proc_21_output_sync_blk[20]);
    assign proc_21_data_FIFO_blk[21] = 1'b0;
    assign proc_21_data_PIPO_blk[21] = 1'b0;
    assign proc_21_start_FIFO_blk[21] = 1'b0;
    assign proc_21_TLF_FIFO_blk[21] = 1'b0;
    assign proc_21_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_21_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_21[21] = dl_detect_out ? proc_dep_vld_vec_21_reg[21] : (proc_21_data_FIFO_blk[21] | proc_21_data_PIPO_blk[21] | proc_21_start_FIFO_blk[21] | proc_21_TLF_FIFO_blk[21] | proc_21_input_sync_blk[21] | proc_21_output_sync_blk[21]);
    assign proc_21_data_FIFO_blk[22] = 1'b0;
    assign proc_21_data_PIPO_blk[22] = 1'b0;
    assign proc_21_start_FIFO_blk[22] = 1'b0;
    assign proc_21_TLF_FIFO_blk[22] = 1'b0;
    assign proc_21_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_21_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_21[22] = dl_detect_out ? proc_dep_vld_vec_21_reg[22] : (proc_21_data_FIFO_blk[22] | proc_21_data_PIPO_blk[22] | proc_21_start_FIFO_blk[22] | proc_21_TLF_FIFO_blk[22] | proc_21_input_sync_blk[22] | proc_21_output_sync_blk[22]);
    assign proc_21_data_FIFO_blk[23] = 1'b0;
    assign proc_21_data_PIPO_blk[23] = 1'b0;
    assign proc_21_start_FIFO_blk[23] = 1'b0;
    assign proc_21_TLF_FIFO_blk[23] = 1'b0;
    assign proc_21_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_21_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_21[23] = dl_detect_out ? proc_dep_vld_vec_21_reg[23] : (proc_21_data_FIFO_blk[23] | proc_21_data_PIPO_blk[23] | proc_21_start_FIFO_blk[23] | proc_21_TLF_FIFO_blk[23] | proc_21_input_sync_blk[23] | proc_21_output_sync_blk[23]);
    assign proc_21_data_FIFO_blk[24] = 1'b0;
    assign proc_21_data_PIPO_blk[24] = 1'b0;
    assign proc_21_start_FIFO_blk[24] = 1'b0;
    assign proc_21_TLF_FIFO_blk[24] = 1'b0;
    assign proc_21_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_21_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_21[24] = dl_detect_out ? proc_dep_vld_vec_21_reg[24] : (proc_21_data_FIFO_blk[24] | proc_21_data_PIPO_blk[24] | proc_21_start_FIFO_blk[24] | proc_21_TLF_FIFO_blk[24] | proc_21_input_sync_blk[24] | proc_21_output_sync_blk[24]);
    assign proc_21_data_FIFO_blk[25] = 1'b0;
    assign proc_21_data_PIPO_blk[25] = 1'b0;
    assign proc_21_start_FIFO_blk[25] = 1'b0;
    assign proc_21_TLF_FIFO_blk[25] = 1'b0;
    assign proc_21_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_21_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_21[25] = dl_detect_out ? proc_dep_vld_vec_21_reg[25] : (proc_21_data_FIFO_blk[25] | proc_21_data_PIPO_blk[25] | proc_21_start_FIFO_blk[25] | proc_21_TLF_FIFO_blk[25] | proc_21_input_sync_blk[25] | proc_21_output_sync_blk[25]);
    assign proc_21_data_FIFO_blk[26] = 1'b0;
    assign proc_21_data_PIPO_blk[26] = 1'b0;
    assign proc_21_start_FIFO_blk[26] = 1'b0;
    assign proc_21_TLF_FIFO_blk[26] = 1'b0;
    assign proc_21_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_21_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_21[26] = dl_detect_out ? proc_dep_vld_vec_21_reg[26] : (proc_21_data_FIFO_blk[26] | proc_21_data_PIPO_blk[26] | proc_21_start_FIFO_blk[26] | proc_21_TLF_FIFO_blk[26] | proc_21_input_sync_blk[26] | proc_21_output_sync_blk[26]);
    assign proc_21_data_FIFO_blk[27] = 1'b0;
    assign proc_21_data_PIPO_blk[27] = 1'b0;
    assign proc_21_start_FIFO_blk[27] = 1'b0;
    assign proc_21_TLF_FIFO_blk[27] = 1'b0;
    assign proc_21_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_21_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_21[27] = dl_detect_out ? proc_dep_vld_vec_21_reg[27] : (proc_21_data_FIFO_blk[27] | proc_21_data_PIPO_blk[27] | proc_21_start_FIFO_blk[27] | proc_21_TLF_FIFO_blk[27] | proc_21_input_sync_blk[27] | proc_21_output_sync_blk[27]);
    assign proc_21_data_FIFO_blk[28] = 1'b0;
    assign proc_21_data_PIPO_blk[28] = 1'b0;
    assign proc_21_start_FIFO_blk[28] = 1'b0;
    assign proc_21_TLF_FIFO_blk[28] = 1'b0;
    assign proc_21_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_21_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_21[28] = dl_detect_out ? proc_dep_vld_vec_21_reg[28] : (proc_21_data_FIFO_blk[28] | proc_21_data_PIPO_blk[28] | proc_21_start_FIFO_blk[28] | proc_21_TLF_FIFO_blk[28] | proc_21_input_sync_blk[28] | proc_21_output_sync_blk[28]);
    assign proc_21_data_FIFO_blk[29] = 1'b0;
    assign proc_21_data_PIPO_blk[29] = 1'b0;
    assign proc_21_start_FIFO_blk[29] = 1'b0;
    assign proc_21_TLF_FIFO_blk[29] = 1'b0;
    assign proc_21_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_21_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_21[29] = dl_detect_out ? proc_dep_vld_vec_21_reg[29] : (proc_21_data_FIFO_blk[29] | proc_21_data_PIPO_blk[29] | proc_21_start_FIFO_blk[29] | proc_21_TLF_FIFO_blk[29] | proc_21_input_sync_blk[29] | proc_21_output_sync_blk[29]);
    assign proc_21_data_FIFO_blk[30] = 1'b0;
    assign proc_21_data_PIPO_blk[30] = 1'b0;
    assign proc_21_start_FIFO_blk[30] = 1'b0;
    assign proc_21_TLF_FIFO_blk[30] = 1'b0;
    assign proc_21_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_21_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_21[30] = dl_detect_out ? proc_dep_vld_vec_21_reg[30] : (proc_21_data_FIFO_blk[30] | proc_21_data_PIPO_blk[30] | proc_21_start_FIFO_blk[30] | proc_21_TLF_FIFO_blk[30] | proc_21_input_sync_blk[30] | proc_21_output_sync_blk[30]);
    assign proc_21_data_FIFO_blk[31] = 1'b0;
    assign proc_21_data_PIPO_blk[31] = 1'b0;
    assign proc_21_start_FIFO_blk[31] = 1'b0;
    assign proc_21_TLF_FIFO_blk[31] = 1'b0;
    assign proc_21_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_21_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_21[31] = dl_detect_out ? proc_dep_vld_vec_21_reg[31] : (proc_21_data_FIFO_blk[31] | proc_21_data_PIPO_blk[31] | proc_21_start_FIFO_blk[31] | proc_21_TLF_FIFO_blk[31] | proc_21_input_sync_blk[31] | proc_21_output_sync_blk[31]);
    assign proc_21_data_FIFO_blk[32] = 1'b0;
    assign proc_21_data_PIPO_blk[32] = 1'b0;
    assign proc_21_start_FIFO_blk[32] = 1'b0;
    assign proc_21_TLF_FIFO_blk[32] = 1'b0;
    assign proc_21_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_16_U0_ap_ready & ProcessingElement_16_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_21_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_21[32] = dl_detect_out ? proc_dep_vld_vec_21_reg[32] : (proc_21_data_FIFO_blk[32] | proc_21_data_PIPO_blk[32] | proc_21_start_FIFO_blk[32] | proc_21_TLF_FIFO_blk[32] | proc_21_input_sync_blk[32] | proc_21_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_21_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_21_reg <= proc_dep_vld_vec_21;
        end
    end
    assign in_chan_dep_vld_vec_21[0] = dep_chan_vld_0_21;
    assign in_chan_dep_data_vec_21[39 : 0] = dep_chan_data_0_21;
    assign token_in_vec_21[0] = token_0_21;
    assign in_chan_dep_vld_vec_21[1] = dep_chan_vld_1_21;
    assign in_chan_dep_data_vec_21[79 : 40] = dep_chan_data_1_21;
    assign token_in_vec_21[1] = token_1_21;
    assign in_chan_dep_vld_vec_21[2] = dep_chan_vld_3_21;
    assign in_chan_dep_data_vec_21[119 : 80] = dep_chan_data_3_21;
    assign token_in_vec_21[2] = token_3_21;
    assign in_chan_dep_vld_vec_21[3] = dep_chan_vld_6_21;
    assign in_chan_dep_data_vec_21[159 : 120] = dep_chan_data_6_21;
    assign token_in_vec_21[3] = token_6_21;
    assign in_chan_dep_vld_vec_21[4] = dep_chan_vld_7_21;
    assign in_chan_dep_data_vec_21[199 : 160] = dep_chan_data_7_21;
    assign token_in_vec_21[4] = token_7_21;
    assign in_chan_dep_vld_vec_21[5] = dep_chan_vld_8_21;
    assign in_chan_dep_data_vec_21[239 : 200] = dep_chan_data_8_21;
    assign token_in_vec_21[5] = token_8_21;
    assign in_chan_dep_vld_vec_21[6] = dep_chan_vld_9_21;
    assign in_chan_dep_data_vec_21[279 : 240] = dep_chan_data_9_21;
    assign token_in_vec_21[6] = token_9_21;
    assign in_chan_dep_vld_vec_21[7] = dep_chan_vld_10_21;
    assign in_chan_dep_data_vec_21[319 : 280] = dep_chan_data_10_21;
    assign token_in_vec_21[7] = token_10_21;
    assign in_chan_dep_vld_vec_21[8] = dep_chan_vld_11_21;
    assign in_chan_dep_data_vec_21[359 : 320] = dep_chan_data_11_21;
    assign token_in_vec_21[8] = token_11_21;
    assign in_chan_dep_vld_vec_21[9] = dep_chan_vld_12_21;
    assign in_chan_dep_data_vec_21[399 : 360] = dep_chan_data_12_21;
    assign token_in_vec_21[9] = token_12_21;
    assign in_chan_dep_vld_vec_21[10] = dep_chan_vld_13_21;
    assign in_chan_dep_data_vec_21[439 : 400] = dep_chan_data_13_21;
    assign token_in_vec_21[10] = token_13_21;
    assign in_chan_dep_vld_vec_21[11] = dep_chan_vld_14_21;
    assign in_chan_dep_data_vec_21[479 : 440] = dep_chan_data_14_21;
    assign token_in_vec_21[11] = token_14_21;
    assign in_chan_dep_vld_vec_21[12] = dep_chan_vld_15_21;
    assign in_chan_dep_data_vec_21[519 : 480] = dep_chan_data_15_21;
    assign token_in_vec_21[12] = token_15_21;
    assign in_chan_dep_vld_vec_21[13] = dep_chan_vld_16_21;
    assign in_chan_dep_data_vec_21[559 : 520] = dep_chan_data_16_21;
    assign token_in_vec_21[13] = token_16_21;
    assign in_chan_dep_vld_vec_21[14] = dep_chan_vld_17_21;
    assign in_chan_dep_data_vec_21[599 : 560] = dep_chan_data_17_21;
    assign token_in_vec_21[14] = token_17_21;
    assign in_chan_dep_vld_vec_21[15] = dep_chan_vld_18_21;
    assign in_chan_dep_data_vec_21[639 : 600] = dep_chan_data_18_21;
    assign token_in_vec_21[15] = token_18_21;
    assign in_chan_dep_vld_vec_21[16] = dep_chan_vld_19_21;
    assign in_chan_dep_data_vec_21[679 : 640] = dep_chan_data_19_21;
    assign token_in_vec_21[16] = token_19_21;
    assign in_chan_dep_vld_vec_21[17] = dep_chan_vld_20_21;
    assign in_chan_dep_data_vec_21[719 : 680] = dep_chan_data_20_21;
    assign token_in_vec_21[17] = token_20_21;
    assign in_chan_dep_vld_vec_21[18] = dep_chan_vld_22_21;
    assign in_chan_dep_data_vec_21[759 : 720] = dep_chan_data_22_21;
    assign token_in_vec_21[18] = token_22_21;
    assign in_chan_dep_vld_vec_21[19] = dep_chan_vld_23_21;
    assign in_chan_dep_data_vec_21[799 : 760] = dep_chan_data_23_21;
    assign token_in_vec_21[19] = token_23_21;
    assign in_chan_dep_vld_vec_21[20] = dep_chan_vld_24_21;
    assign in_chan_dep_data_vec_21[839 : 800] = dep_chan_data_24_21;
    assign token_in_vec_21[20] = token_24_21;
    assign in_chan_dep_vld_vec_21[21] = dep_chan_vld_25_21;
    assign in_chan_dep_data_vec_21[879 : 840] = dep_chan_data_25_21;
    assign token_in_vec_21[21] = token_25_21;
    assign in_chan_dep_vld_vec_21[22] = dep_chan_vld_26_21;
    assign in_chan_dep_data_vec_21[919 : 880] = dep_chan_data_26_21;
    assign token_in_vec_21[22] = token_26_21;
    assign in_chan_dep_vld_vec_21[23] = dep_chan_vld_27_21;
    assign in_chan_dep_data_vec_21[959 : 920] = dep_chan_data_27_21;
    assign token_in_vec_21[23] = token_27_21;
    assign in_chan_dep_vld_vec_21[24] = dep_chan_vld_28_21;
    assign in_chan_dep_data_vec_21[999 : 960] = dep_chan_data_28_21;
    assign token_in_vec_21[24] = token_28_21;
    assign in_chan_dep_vld_vec_21[25] = dep_chan_vld_29_21;
    assign in_chan_dep_data_vec_21[1039 : 1000] = dep_chan_data_29_21;
    assign token_in_vec_21[25] = token_29_21;
    assign in_chan_dep_vld_vec_21[26] = dep_chan_vld_30_21;
    assign in_chan_dep_data_vec_21[1079 : 1040] = dep_chan_data_30_21;
    assign token_in_vec_21[26] = token_30_21;
    assign in_chan_dep_vld_vec_21[27] = dep_chan_vld_31_21;
    assign in_chan_dep_data_vec_21[1119 : 1080] = dep_chan_data_31_21;
    assign token_in_vec_21[27] = token_31_21;
    assign in_chan_dep_vld_vec_21[28] = dep_chan_vld_32_21;
    assign in_chan_dep_data_vec_21[1159 : 1120] = dep_chan_data_32_21;
    assign token_in_vec_21[28] = token_32_21;
    assign in_chan_dep_vld_vec_21[29] = dep_chan_vld_33_21;
    assign in_chan_dep_data_vec_21[1199 : 1160] = dep_chan_data_33_21;
    assign token_in_vec_21[29] = token_33_21;
    assign in_chan_dep_vld_vec_21[30] = dep_chan_vld_34_21;
    assign in_chan_dep_data_vec_21[1239 : 1200] = dep_chan_data_34_21;
    assign token_in_vec_21[30] = token_34_21;
    assign in_chan_dep_vld_vec_21[31] = dep_chan_vld_35_21;
    assign in_chan_dep_data_vec_21[1279 : 1240] = dep_chan_data_35_21;
    assign token_in_vec_21[31] = token_35_21;
    assign in_chan_dep_vld_vec_21[32] = dep_chan_vld_36_21;
    assign in_chan_dep_data_vec_21[1319 : 1280] = dep_chan_data_36_21;
    assign token_in_vec_21[32] = token_36_21;
    assign dep_chan_vld_21_20 = out_chan_dep_vld_vec_21[0];
    assign dep_chan_data_21_20 = out_chan_dep_data_21;
    assign token_21_20 = token_out_vec_21[0];
    assign dep_chan_vld_21_22 = out_chan_dep_vld_vec_21[1];
    assign dep_chan_data_21_22 = out_chan_dep_data_21;
    assign token_21_22 = token_out_vec_21[1];
    assign dep_chan_vld_21_0 = out_chan_dep_vld_vec_21[2];
    assign dep_chan_data_21_0 = out_chan_dep_data_21;
    assign token_21_0 = token_out_vec_21[2];
    assign dep_chan_vld_21_1 = out_chan_dep_vld_vec_21[3];
    assign dep_chan_data_21_1 = out_chan_dep_data_21;
    assign token_21_1 = token_out_vec_21[3];
    assign dep_chan_vld_21_3 = out_chan_dep_vld_vec_21[4];
    assign dep_chan_data_21_3 = out_chan_dep_data_21;
    assign token_21_3 = token_out_vec_21[4];
    assign dep_chan_vld_21_6 = out_chan_dep_vld_vec_21[5];
    assign dep_chan_data_21_6 = out_chan_dep_data_21;
    assign token_21_6 = token_out_vec_21[5];
    assign dep_chan_vld_21_7 = out_chan_dep_vld_vec_21[6];
    assign dep_chan_data_21_7 = out_chan_dep_data_21;
    assign token_21_7 = token_out_vec_21[6];
    assign dep_chan_vld_21_8 = out_chan_dep_vld_vec_21[7];
    assign dep_chan_data_21_8 = out_chan_dep_data_21;
    assign token_21_8 = token_out_vec_21[7];
    assign dep_chan_vld_21_9 = out_chan_dep_vld_vec_21[8];
    assign dep_chan_data_21_9 = out_chan_dep_data_21;
    assign token_21_9 = token_out_vec_21[8];
    assign dep_chan_vld_21_10 = out_chan_dep_vld_vec_21[9];
    assign dep_chan_data_21_10 = out_chan_dep_data_21;
    assign token_21_10 = token_out_vec_21[9];
    assign dep_chan_vld_21_11 = out_chan_dep_vld_vec_21[10];
    assign dep_chan_data_21_11 = out_chan_dep_data_21;
    assign token_21_11 = token_out_vec_21[10];
    assign dep_chan_vld_21_12 = out_chan_dep_vld_vec_21[11];
    assign dep_chan_data_21_12 = out_chan_dep_data_21;
    assign token_21_12 = token_out_vec_21[11];
    assign dep_chan_vld_21_13 = out_chan_dep_vld_vec_21[12];
    assign dep_chan_data_21_13 = out_chan_dep_data_21;
    assign token_21_13 = token_out_vec_21[12];
    assign dep_chan_vld_21_14 = out_chan_dep_vld_vec_21[13];
    assign dep_chan_data_21_14 = out_chan_dep_data_21;
    assign token_21_14 = token_out_vec_21[13];
    assign dep_chan_vld_21_15 = out_chan_dep_vld_vec_21[14];
    assign dep_chan_data_21_15 = out_chan_dep_data_21;
    assign token_21_15 = token_out_vec_21[14];
    assign dep_chan_vld_21_16 = out_chan_dep_vld_vec_21[15];
    assign dep_chan_data_21_16 = out_chan_dep_data_21;
    assign token_21_16 = token_out_vec_21[15];
    assign dep_chan_vld_21_17 = out_chan_dep_vld_vec_21[16];
    assign dep_chan_data_21_17 = out_chan_dep_data_21;
    assign token_21_17 = token_out_vec_21[16];
    assign dep_chan_vld_21_18 = out_chan_dep_vld_vec_21[17];
    assign dep_chan_data_21_18 = out_chan_dep_data_21;
    assign token_21_18 = token_out_vec_21[17];
    assign dep_chan_vld_21_19 = out_chan_dep_vld_vec_21[18];
    assign dep_chan_data_21_19 = out_chan_dep_data_21;
    assign token_21_19 = token_out_vec_21[18];
    assign dep_chan_vld_21_23 = out_chan_dep_vld_vec_21[19];
    assign dep_chan_data_21_23 = out_chan_dep_data_21;
    assign token_21_23 = token_out_vec_21[19];
    assign dep_chan_vld_21_24 = out_chan_dep_vld_vec_21[20];
    assign dep_chan_data_21_24 = out_chan_dep_data_21;
    assign token_21_24 = token_out_vec_21[20];
    assign dep_chan_vld_21_25 = out_chan_dep_vld_vec_21[21];
    assign dep_chan_data_21_25 = out_chan_dep_data_21;
    assign token_21_25 = token_out_vec_21[21];
    assign dep_chan_vld_21_26 = out_chan_dep_vld_vec_21[22];
    assign dep_chan_data_21_26 = out_chan_dep_data_21;
    assign token_21_26 = token_out_vec_21[22];
    assign dep_chan_vld_21_27 = out_chan_dep_vld_vec_21[23];
    assign dep_chan_data_21_27 = out_chan_dep_data_21;
    assign token_21_27 = token_out_vec_21[23];
    assign dep_chan_vld_21_28 = out_chan_dep_vld_vec_21[24];
    assign dep_chan_data_21_28 = out_chan_dep_data_21;
    assign token_21_28 = token_out_vec_21[24];
    assign dep_chan_vld_21_29 = out_chan_dep_vld_vec_21[25];
    assign dep_chan_data_21_29 = out_chan_dep_data_21;
    assign token_21_29 = token_out_vec_21[25];
    assign dep_chan_vld_21_30 = out_chan_dep_vld_vec_21[26];
    assign dep_chan_data_21_30 = out_chan_dep_data_21;
    assign token_21_30 = token_out_vec_21[26];
    assign dep_chan_vld_21_31 = out_chan_dep_vld_vec_21[27];
    assign dep_chan_data_21_31 = out_chan_dep_data_21;
    assign token_21_31 = token_out_vec_21[27];
    assign dep_chan_vld_21_32 = out_chan_dep_vld_vec_21[28];
    assign dep_chan_data_21_32 = out_chan_dep_data_21;
    assign token_21_32 = token_out_vec_21[28];
    assign dep_chan_vld_21_33 = out_chan_dep_vld_vec_21[29];
    assign dep_chan_data_21_33 = out_chan_dep_data_21;
    assign token_21_33 = token_out_vec_21[29];
    assign dep_chan_vld_21_34 = out_chan_dep_vld_vec_21[30];
    assign dep_chan_data_21_34 = out_chan_dep_data_21;
    assign token_21_34 = token_out_vec_21[30];
    assign dep_chan_vld_21_35 = out_chan_dep_vld_vec_21[31];
    assign dep_chan_data_21_35 = out_chan_dep_data_21;
    assign token_21_35 = token_out_vec_21[31];
    assign dep_chan_vld_21_36 = out_chan_dep_vld_vec_21[32];
    assign dep_chan_data_21_36 = out_chan_dep_data_21;
    assign token_21_36 = token_out_vec_21[32];

    // Process: ProcessingElement_17_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 22, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_22 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_22),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_22),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_22),
        .token_in_vec(token_in_vec_22),
        .dl_detect_in(dl_detect_out),
        .origin(origin[22]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_22),
        .out_chan_dep_data(out_chan_dep_data_22),
        .token_out_vec(token_out_vec_22),
        .dl_detect_out(dl_in_vec[22]));

    assign proc_22_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_16_blk_n) | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_16_blk_n) | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_WriteC_Flattened_fu_179.cPipes_16_blk_n);
    assign proc_22_data_PIPO_blk[0] = 1'b0;
    assign proc_22_start_FIFO_blk[0] = 1'b0;
    assign proc_22_TLF_FIFO_blk[0] = 1'b0;
    assign proc_22_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_22_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_22[0] = dl_detect_out ? proc_dep_vld_vec_22_reg[0] : (proc_22_data_FIFO_blk[0] | proc_22_data_PIPO_blk[0] | proc_22_start_FIFO_blk[0] | proc_22_TLF_FIFO_blk[0] | proc_22_input_sync_blk[0] | proc_22_output_sync_blk[0]);
    assign proc_22_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_17_blk_n) | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_17_blk_n) | (~ProcessingElement_17_U0.grp_ProcessingElement_17_Pipeline_WriteC_Flattened_fu_179.cPipes_17_blk_n);
    assign proc_22_data_PIPO_blk[1] = 1'b0;
    assign proc_22_start_FIFO_blk[1] = 1'b0;
    assign proc_22_TLF_FIFO_blk[1] = 1'b0;
    assign proc_22_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_22_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_22[1] = dl_detect_out ? proc_dep_vld_vec_22_reg[1] : (proc_22_data_FIFO_blk[1] | proc_22_data_PIPO_blk[1] | proc_22_start_FIFO_blk[1] | proc_22_TLF_FIFO_blk[1] | proc_22_input_sync_blk[1] | proc_22_output_sync_blk[1]);
    assign proc_22_data_FIFO_blk[2] = 1'b0;
    assign proc_22_data_PIPO_blk[2] = 1'b0;
    assign proc_22_start_FIFO_blk[2] = 1'b0;
    assign proc_22_TLF_FIFO_blk[2] = 1'b0;
    assign proc_22_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_22_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_22[2] = dl_detect_out ? proc_dep_vld_vec_22_reg[2] : (proc_22_data_FIFO_blk[2] | proc_22_data_PIPO_blk[2] | proc_22_start_FIFO_blk[2] | proc_22_TLF_FIFO_blk[2] | proc_22_input_sync_blk[2] | proc_22_output_sync_blk[2]);
    assign proc_22_data_FIFO_blk[3] = 1'b0;
    assign proc_22_data_PIPO_blk[3] = 1'b0;
    assign proc_22_start_FIFO_blk[3] = 1'b0;
    assign proc_22_TLF_FIFO_blk[3] = 1'b0;
    assign proc_22_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_22_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_22[3] = dl_detect_out ? proc_dep_vld_vec_22_reg[3] : (proc_22_data_FIFO_blk[3] | proc_22_data_PIPO_blk[3] | proc_22_start_FIFO_blk[3] | proc_22_TLF_FIFO_blk[3] | proc_22_input_sync_blk[3] | proc_22_output_sync_blk[3]);
    assign proc_22_data_FIFO_blk[4] = 1'b0;
    assign proc_22_data_PIPO_blk[4] = 1'b0;
    assign proc_22_start_FIFO_blk[4] = 1'b0;
    assign proc_22_TLF_FIFO_blk[4] = 1'b0;
    assign proc_22_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_22_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_22[4] = dl_detect_out ? proc_dep_vld_vec_22_reg[4] : (proc_22_data_FIFO_blk[4] | proc_22_data_PIPO_blk[4] | proc_22_start_FIFO_blk[4] | proc_22_TLF_FIFO_blk[4] | proc_22_input_sync_blk[4] | proc_22_output_sync_blk[4]);
    assign proc_22_data_FIFO_blk[5] = 1'b0;
    assign proc_22_data_PIPO_blk[5] = 1'b0;
    assign proc_22_start_FIFO_blk[5] = 1'b0;
    assign proc_22_TLF_FIFO_blk[5] = 1'b0;
    assign proc_22_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_22_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_22[5] = dl_detect_out ? proc_dep_vld_vec_22_reg[5] : (proc_22_data_FIFO_blk[5] | proc_22_data_PIPO_blk[5] | proc_22_start_FIFO_blk[5] | proc_22_TLF_FIFO_blk[5] | proc_22_input_sync_blk[5] | proc_22_output_sync_blk[5]);
    assign proc_22_data_FIFO_blk[6] = 1'b0;
    assign proc_22_data_PIPO_blk[6] = 1'b0;
    assign proc_22_start_FIFO_blk[6] = 1'b0;
    assign proc_22_TLF_FIFO_blk[6] = 1'b0;
    assign proc_22_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_22_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_22[6] = dl_detect_out ? proc_dep_vld_vec_22_reg[6] : (proc_22_data_FIFO_blk[6] | proc_22_data_PIPO_blk[6] | proc_22_start_FIFO_blk[6] | proc_22_TLF_FIFO_blk[6] | proc_22_input_sync_blk[6] | proc_22_output_sync_blk[6]);
    assign proc_22_data_FIFO_blk[7] = 1'b0;
    assign proc_22_data_PIPO_blk[7] = 1'b0;
    assign proc_22_start_FIFO_blk[7] = 1'b0;
    assign proc_22_TLF_FIFO_blk[7] = 1'b0;
    assign proc_22_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_22_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_22[7] = dl_detect_out ? proc_dep_vld_vec_22_reg[7] : (proc_22_data_FIFO_blk[7] | proc_22_data_PIPO_blk[7] | proc_22_start_FIFO_blk[7] | proc_22_TLF_FIFO_blk[7] | proc_22_input_sync_blk[7] | proc_22_output_sync_blk[7]);
    assign proc_22_data_FIFO_blk[8] = 1'b0;
    assign proc_22_data_PIPO_blk[8] = 1'b0;
    assign proc_22_start_FIFO_blk[8] = 1'b0;
    assign proc_22_TLF_FIFO_blk[8] = 1'b0;
    assign proc_22_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_22_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_22[8] = dl_detect_out ? proc_dep_vld_vec_22_reg[8] : (proc_22_data_FIFO_blk[8] | proc_22_data_PIPO_blk[8] | proc_22_start_FIFO_blk[8] | proc_22_TLF_FIFO_blk[8] | proc_22_input_sync_blk[8] | proc_22_output_sync_blk[8]);
    assign proc_22_data_FIFO_blk[9] = 1'b0;
    assign proc_22_data_PIPO_blk[9] = 1'b0;
    assign proc_22_start_FIFO_blk[9] = 1'b0;
    assign proc_22_TLF_FIFO_blk[9] = 1'b0;
    assign proc_22_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_22_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_22[9] = dl_detect_out ? proc_dep_vld_vec_22_reg[9] : (proc_22_data_FIFO_blk[9] | proc_22_data_PIPO_blk[9] | proc_22_start_FIFO_blk[9] | proc_22_TLF_FIFO_blk[9] | proc_22_input_sync_blk[9] | proc_22_output_sync_blk[9]);
    assign proc_22_data_FIFO_blk[10] = 1'b0;
    assign proc_22_data_PIPO_blk[10] = 1'b0;
    assign proc_22_start_FIFO_blk[10] = 1'b0;
    assign proc_22_TLF_FIFO_blk[10] = 1'b0;
    assign proc_22_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_22_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_22[10] = dl_detect_out ? proc_dep_vld_vec_22_reg[10] : (proc_22_data_FIFO_blk[10] | proc_22_data_PIPO_blk[10] | proc_22_start_FIFO_blk[10] | proc_22_TLF_FIFO_blk[10] | proc_22_input_sync_blk[10] | proc_22_output_sync_blk[10]);
    assign proc_22_data_FIFO_blk[11] = 1'b0;
    assign proc_22_data_PIPO_blk[11] = 1'b0;
    assign proc_22_start_FIFO_blk[11] = 1'b0;
    assign proc_22_TLF_FIFO_blk[11] = 1'b0;
    assign proc_22_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_22_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_22[11] = dl_detect_out ? proc_dep_vld_vec_22_reg[11] : (proc_22_data_FIFO_blk[11] | proc_22_data_PIPO_blk[11] | proc_22_start_FIFO_blk[11] | proc_22_TLF_FIFO_blk[11] | proc_22_input_sync_blk[11] | proc_22_output_sync_blk[11]);
    assign proc_22_data_FIFO_blk[12] = 1'b0;
    assign proc_22_data_PIPO_blk[12] = 1'b0;
    assign proc_22_start_FIFO_blk[12] = 1'b0;
    assign proc_22_TLF_FIFO_blk[12] = 1'b0;
    assign proc_22_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_22_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_22[12] = dl_detect_out ? proc_dep_vld_vec_22_reg[12] : (proc_22_data_FIFO_blk[12] | proc_22_data_PIPO_blk[12] | proc_22_start_FIFO_blk[12] | proc_22_TLF_FIFO_blk[12] | proc_22_input_sync_blk[12] | proc_22_output_sync_blk[12]);
    assign proc_22_data_FIFO_blk[13] = 1'b0;
    assign proc_22_data_PIPO_blk[13] = 1'b0;
    assign proc_22_start_FIFO_blk[13] = 1'b0;
    assign proc_22_TLF_FIFO_blk[13] = 1'b0;
    assign proc_22_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_22_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_22[13] = dl_detect_out ? proc_dep_vld_vec_22_reg[13] : (proc_22_data_FIFO_blk[13] | proc_22_data_PIPO_blk[13] | proc_22_start_FIFO_blk[13] | proc_22_TLF_FIFO_blk[13] | proc_22_input_sync_blk[13] | proc_22_output_sync_blk[13]);
    assign proc_22_data_FIFO_blk[14] = 1'b0;
    assign proc_22_data_PIPO_blk[14] = 1'b0;
    assign proc_22_start_FIFO_blk[14] = 1'b0;
    assign proc_22_TLF_FIFO_blk[14] = 1'b0;
    assign proc_22_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_22_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_22[14] = dl_detect_out ? proc_dep_vld_vec_22_reg[14] : (proc_22_data_FIFO_blk[14] | proc_22_data_PIPO_blk[14] | proc_22_start_FIFO_blk[14] | proc_22_TLF_FIFO_blk[14] | proc_22_input_sync_blk[14] | proc_22_output_sync_blk[14]);
    assign proc_22_data_FIFO_blk[15] = 1'b0;
    assign proc_22_data_PIPO_blk[15] = 1'b0;
    assign proc_22_start_FIFO_blk[15] = 1'b0;
    assign proc_22_TLF_FIFO_blk[15] = 1'b0;
    assign proc_22_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_22_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_22[15] = dl_detect_out ? proc_dep_vld_vec_22_reg[15] : (proc_22_data_FIFO_blk[15] | proc_22_data_PIPO_blk[15] | proc_22_start_FIFO_blk[15] | proc_22_TLF_FIFO_blk[15] | proc_22_input_sync_blk[15] | proc_22_output_sync_blk[15]);
    assign proc_22_data_FIFO_blk[16] = 1'b0;
    assign proc_22_data_PIPO_blk[16] = 1'b0;
    assign proc_22_start_FIFO_blk[16] = 1'b0;
    assign proc_22_TLF_FIFO_blk[16] = 1'b0;
    assign proc_22_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_22_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_22[16] = dl_detect_out ? proc_dep_vld_vec_22_reg[16] : (proc_22_data_FIFO_blk[16] | proc_22_data_PIPO_blk[16] | proc_22_start_FIFO_blk[16] | proc_22_TLF_FIFO_blk[16] | proc_22_input_sync_blk[16] | proc_22_output_sync_blk[16]);
    assign proc_22_data_FIFO_blk[17] = 1'b0;
    assign proc_22_data_PIPO_blk[17] = 1'b0;
    assign proc_22_start_FIFO_blk[17] = 1'b0;
    assign proc_22_TLF_FIFO_blk[17] = 1'b0;
    assign proc_22_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_22_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_22[17] = dl_detect_out ? proc_dep_vld_vec_22_reg[17] : (proc_22_data_FIFO_blk[17] | proc_22_data_PIPO_blk[17] | proc_22_start_FIFO_blk[17] | proc_22_TLF_FIFO_blk[17] | proc_22_input_sync_blk[17] | proc_22_output_sync_blk[17]);
    assign proc_22_data_FIFO_blk[18] = 1'b0;
    assign proc_22_data_PIPO_blk[18] = 1'b0;
    assign proc_22_start_FIFO_blk[18] = 1'b0;
    assign proc_22_TLF_FIFO_blk[18] = 1'b0;
    assign proc_22_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_22_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_22[18] = dl_detect_out ? proc_dep_vld_vec_22_reg[18] : (proc_22_data_FIFO_blk[18] | proc_22_data_PIPO_blk[18] | proc_22_start_FIFO_blk[18] | proc_22_TLF_FIFO_blk[18] | proc_22_input_sync_blk[18] | proc_22_output_sync_blk[18]);
    assign proc_22_data_FIFO_blk[19] = 1'b0;
    assign proc_22_data_PIPO_blk[19] = 1'b0;
    assign proc_22_start_FIFO_blk[19] = 1'b0;
    assign proc_22_TLF_FIFO_blk[19] = 1'b0;
    assign proc_22_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_22_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_22[19] = dl_detect_out ? proc_dep_vld_vec_22_reg[19] : (proc_22_data_FIFO_blk[19] | proc_22_data_PIPO_blk[19] | proc_22_start_FIFO_blk[19] | proc_22_TLF_FIFO_blk[19] | proc_22_input_sync_blk[19] | proc_22_output_sync_blk[19]);
    assign proc_22_data_FIFO_blk[20] = 1'b0;
    assign proc_22_data_PIPO_blk[20] = 1'b0;
    assign proc_22_start_FIFO_blk[20] = 1'b0;
    assign proc_22_TLF_FIFO_blk[20] = 1'b0;
    assign proc_22_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_22_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_22[20] = dl_detect_out ? proc_dep_vld_vec_22_reg[20] : (proc_22_data_FIFO_blk[20] | proc_22_data_PIPO_blk[20] | proc_22_start_FIFO_blk[20] | proc_22_TLF_FIFO_blk[20] | proc_22_input_sync_blk[20] | proc_22_output_sync_blk[20]);
    assign proc_22_data_FIFO_blk[21] = 1'b0;
    assign proc_22_data_PIPO_blk[21] = 1'b0;
    assign proc_22_start_FIFO_blk[21] = 1'b0;
    assign proc_22_TLF_FIFO_blk[21] = 1'b0;
    assign proc_22_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_22_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_22[21] = dl_detect_out ? proc_dep_vld_vec_22_reg[21] : (proc_22_data_FIFO_blk[21] | proc_22_data_PIPO_blk[21] | proc_22_start_FIFO_blk[21] | proc_22_TLF_FIFO_blk[21] | proc_22_input_sync_blk[21] | proc_22_output_sync_blk[21]);
    assign proc_22_data_FIFO_blk[22] = 1'b0;
    assign proc_22_data_PIPO_blk[22] = 1'b0;
    assign proc_22_start_FIFO_blk[22] = 1'b0;
    assign proc_22_TLF_FIFO_blk[22] = 1'b0;
    assign proc_22_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_22_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_22[22] = dl_detect_out ? proc_dep_vld_vec_22_reg[22] : (proc_22_data_FIFO_blk[22] | proc_22_data_PIPO_blk[22] | proc_22_start_FIFO_blk[22] | proc_22_TLF_FIFO_blk[22] | proc_22_input_sync_blk[22] | proc_22_output_sync_blk[22]);
    assign proc_22_data_FIFO_blk[23] = 1'b0;
    assign proc_22_data_PIPO_blk[23] = 1'b0;
    assign proc_22_start_FIFO_blk[23] = 1'b0;
    assign proc_22_TLF_FIFO_blk[23] = 1'b0;
    assign proc_22_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_22_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_22[23] = dl_detect_out ? proc_dep_vld_vec_22_reg[23] : (proc_22_data_FIFO_blk[23] | proc_22_data_PIPO_blk[23] | proc_22_start_FIFO_blk[23] | proc_22_TLF_FIFO_blk[23] | proc_22_input_sync_blk[23] | proc_22_output_sync_blk[23]);
    assign proc_22_data_FIFO_blk[24] = 1'b0;
    assign proc_22_data_PIPO_blk[24] = 1'b0;
    assign proc_22_start_FIFO_blk[24] = 1'b0;
    assign proc_22_TLF_FIFO_blk[24] = 1'b0;
    assign proc_22_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_22_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_22[24] = dl_detect_out ? proc_dep_vld_vec_22_reg[24] : (proc_22_data_FIFO_blk[24] | proc_22_data_PIPO_blk[24] | proc_22_start_FIFO_blk[24] | proc_22_TLF_FIFO_blk[24] | proc_22_input_sync_blk[24] | proc_22_output_sync_blk[24]);
    assign proc_22_data_FIFO_blk[25] = 1'b0;
    assign proc_22_data_PIPO_blk[25] = 1'b0;
    assign proc_22_start_FIFO_blk[25] = 1'b0;
    assign proc_22_TLF_FIFO_blk[25] = 1'b0;
    assign proc_22_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_22_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_22[25] = dl_detect_out ? proc_dep_vld_vec_22_reg[25] : (proc_22_data_FIFO_blk[25] | proc_22_data_PIPO_blk[25] | proc_22_start_FIFO_blk[25] | proc_22_TLF_FIFO_blk[25] | proc_22_input_sync_blk[25] | proc_22_output_sync_blk[25]);
    assign proc_22_data_FIFO_blk[26] = 1'b0;
    assign proc_22_data_PIPO_blk[26] = 1'b0;
    assign proc_22_start_FIFO_blk[26] = 1'b0;
    assign proc_22_TLF_FIFO_blk[26] = 1'b0;
    assign proc_22_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_22_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_22[26] = dl_detect_out ? proc_dep_vld_vec_22_reg[26] : (proc_22_data_FIFO_blk[26] | proc_22_data_PIPO_blk[26] | proc_22_start_FIFO_blk[26] | proc_22_TLF_FIFO_blk[26] | proc_22_input_sync_blk[26] | proc_22_output_sync_blk[26]);
    assign proc_22_data_FIFO_blk[27] = 1'b0;
    assign proc_22_data_PIPO_blk[27] = 1'b0;
    assign proc_22_start_FIFO_blk[27] = 1'b0;
    assign proc_22_TLF_FIFO_blk[27] = 1'b0;
    assign proc_22_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_22_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_22[27] = dl_detect_out ? proc_dep_vld_vec_22_reg[27] : (proc_22_data_FIFO_blk[27] | proc_22_data_PIPO_blk[27] | proc_22_start_FIFO_blk[27] | proc_22_TLF_FIFO_blk[27] | proc_22_input_sync_blk[27] | proc_22_output_sync_blk[27]);
    assign proc_22_data_FIFO_blk[28] = 1'b0;
    assign proc_22_data_PIPO_blk[28] = 1'b0;
    assign proc_22_start_FIFO_blk[28] = 1'b0;
    assign proc_22_TLF_FIFO_blk[28] = 1'b0;
    assign proc_22_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_22_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_22[28] = dl_detect_out ? proc_dep_vld_vec_22_reg[28] : (proc_22_data_FIFO_blk[28] | proc_22_data_PIPO_blk[28] | proc_22_start_FIFO_blk[28] | proc_22_TLF_FIFO_blk[28] | proc_22_input_sync_blk[28] | proc_22_output_sync_blk[28]);
    assign proc_22_data_FIFO_blk[29] = 1'b0;
    assign proc_22_data_PIPO_blk[29] = 1'b0;
    assign proc_22_start_FIFO_blk[29] = 1'b0;
    assign proc_22_TLF_FIFO_blk[29] = 1'b0;
    assign proc_22_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_22_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_22[29] = dl_detect_out ? proc_dep_vld_vec_22_reg[29] : (proc_22_data_FIFO_blk[29] | proc_22_data_PIPO_blk[29] | proc_22_start_FIFO_blk[29] | proc_22_TLF_FIFO_blk[29] | proc_22_input_sync_blk[29] | proc_22_output_sync_blk[29]);
    assign proc_22_data_FIFO_blk[30] = 1'b0;
    assign proc_22_data_PIPO_blk[30] = 1'b0;
    assign proc_22_start_FIFO_blk[30] = 1'b0;
    assign proc_22_TLF_FIFO_blk[30] = 1'b0;
    assign proc_22_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_22_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_22[30] = dl_detect_out ? proc_dep_vld_vec_22_reg[30] : (proc_22_data_FIFO_blk[30] | proc_22_data_PIPO_blk[30] | proc_22_start_FIFO_blk[30] | proc_22_TLF_FIFO_blk[30] | proc_22_input_sync_blk[30] | proc_22_output_sync_blk[30]);
    assign proc_22_data_FIFO_blk[31] = 1'b0;
    assign proc_22_data_PIPO_blk[31] = 1'b0;
    assign proc_22_start_FIFO_blk[31] = 1'b0;
    assign proc_22_TLF_FIFO_blk[31] = 1'b0;
    assign proc_22_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_22_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_22[31] = dl_detect_out ? proc_dep_vld_vec_22_reg[31] : (proc_22_data_FIFO_blk[31] | proc_22_data_PIPO_blk[31] | proc_22_start_FIFO_blk[31] | proc_22_TLF_FIFO_blk[31] | proc_22_input_sync_blk[31] | proc_22_output_sync_blk[31]);
    assign proc_22_data_FIFO_blk[32] = 1'b0;
    assign proc_22_data_PIPO_blk[32] = 1'b0;
    assign proc_22_start_FIFO_blk[32] = 1'b0;
    assign proc_22_TLF_FIFO_blk[32] = 1'b0;
    assign proc_22_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_17_U0_ap_ready & ProcessingElement_17_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_22_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_22[32] = dl_detect_out ? proc_dep_vld_vec_22_reg[32] : (proc_22_data_FIFO_blk[32] | proc_22_data_PIPO_blk[32] | proc_22_start_FIFO_blk[32] | proc_22_TLF_FIFO_blk[32] | proc_22_input_sync_blk[32] | proc_22_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_22_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_22_reg <= proc_dep_vld_vec_22;
        end
    end
    assign in_chan_dep_vld_vec_22[0] = dep_chan_vld_0_22;
    assign in_chan_dep_data_vec_22[39 : 0] = dep_chan_data_0_22;
    assign token_in_vec_22[0] = token_0_22;
    assign in_chan_dep_vld_vec_22[1] = dep_chan_vld_1_22;
    assign in_chan_dep_data_vec_22[79 : 40] = dep_chan_data_1_22;
    assign token_in_vec_22[1] = token_1_22;
    assign in_chan_dep_vld_vec_22[2] = dep_chan_vld_3_22;
    assign in_chan_dep_data_vec_22[119 : 80] = dep_chan_data_3_22;
    assign token_in_vec_22[2] = token_3_22;
    assign in_chan_dep_vld_vec_22[3] = dep_chan_vld_6_22;
    assign in_chan_dep_data_vec_22[159 : 120] = dep_chan_data_6_22;
    assign token_in_vec_22[3] = token_6_22;
    assign in_chan_dep_vld_vec_22[4] = dep_chan_vld_7_22;
    assign in_chan_dep_data_vec_22[199 : 160] = dep_chan_data_7_22;
    assign token_in_vec_22[4] = token_7_22;
    assign in_chan_dep_vld_vec_22[5] = dep_chan_vld_8_22;
    assign in_chan_dep_data_vec_22[239 : 200] = dep_chan_data_8_22;
    assign token_in_vec_22[5] = token_8_22;
    assign in_chan_dep_vld_vec_22[6] = dep_chan_vld_9_22;
    assign in_chan_dep_data_vec_22[279 : 240] = dep_chan_data_9_22;
    assign token_in_vec_22[6] = token_9_22;
    assign in_chan_dep_vld_vec_22[7] = dep_chan_vld_10_22;
    assign in_chan_dep_data_vec_22[319 : 280] = dep_chan_data_10_22;
    assign token_in_vec_22[7] = token_10_22;
    assign in_chan_dep_vld_vec_22[8] = dep_chan_vld_11_22;
    assign in_chan_dep_data_vec_22[359 : 320] = dep_chan_data_11_22;
    assign token_in_vec_22[8] = token_11_22;
    assign in_chan_dep_vld_vec_22[9] = dep_chan_vld_12_22;
    assign in_chan_dep_data_vec_22[399 : 360] = dep_chan_data_12_22;
    assign token_in_vec_22[9] = token_12_22;
    assign in_chan_dep_vld_vec_22[10] = dep_chan_vld_13_22;
    assign in_chan_dep_data_vec_22[439 : 400] = dep_chan_data_13_22;
    assign token_in_vec_22[10] = token_13_22;
    assign in_chan_dep_vld_vec_22[11] = dep_chan_vld_14_22;
    assign in_chan_dep_data_vec_22[479 : 440] = dep_chan_data_14_22;
    assign token_in_vec_22[11] = token_14_22;
    assign in_chan_dep_vld_vec_22[12] = dep_chan_vld_15_22;
    assign in_chan_dep_data_vec_22[519 : 480] = dep_chan_data_15_22;
    assign token_in_vec_22[12] = token_15_22;
    assign in_chan_dep_vld_vec_22[13] = dep_chan_vld_16_22;
    assign in_chan_dep_data_vec_22[559 : 520] = dep_chan_data_16_22;
    assign token_in_vec_22[13] = token_16_22;
    assign in_chan_dep_vld_vec_22[14] = dep_chan_vld_17_22;
    assign in_chan_dep_data_vec_22[599 : 560] = dep_chan_data_17_22;
    assign token_in_vec_22[14] = token_17_22;
    assign in_chan_dep_vld_vec_22[15] = dep_chan_vld_18_22;
    assign in_chan_dep_data_vec_22[639 : 600] = dep_chan_data_18_22;
    assign token_in_vec_22[15] = token_18_22;
    assign in_chan_dep_vld_vec_22[16] = dep_chan_vld_19_22;
    assign in_chan_dep_data_vec_22[679 : 640] = dep_chan_data_19_22;
    assign token_in_vec_22[16] = token_19_22;
    assign in_chan_dep_vld_vec_22[17] = dep_chan_vld_20_22;
    assign in_chan_dep_data_vec_22[719 : 680] = dep_chan_data_20_22;
    assign token_in_vec_22[17] = token_20_22;
    assign in_chan_dep_vld_vec_22[18] = dep_chan_vld_21_22;
    assign in_chan_dep_data_vec_22[759 : 720] = dep_chan_data_21_22;
    assign token_in_vec_22[18] = token_21_22;
    assign in_chan_dep_vld_vec_22[19] = dep_chan_vld_23_22;
    assign in_chan_dep_data_vec_22[799 : 760] = dep_chan_data_23_22;
    assign token_in_vec_22[19] = token_23_22;
    assign in_chan_dep_vld_vec_22[20] = dep_chan_vld_24_22;
    assign in_chan_dep_data_vec_22[839 : 800] = dep_chan_data_24_22;
    assign token_in_vec_22[20] = token_24_22;
    assign in_chan_dep_vld_vec_22[21] = dep_chan_vld_25_22;
    assign in_chan_dep_data_vec_22[879 : 840] = dep_chan_data_25_22;
    assign token_in_vec_22[21] = token_25_22;
    assign in_chan_dep_vld_vec_22[22] = dep_chan_vld_26_22;
    assign in_chan_dep_data_vec_22[919 : 880] = dep_chan_data_26_22;
    assign token_in_vec_22[22] = token_26_22;
    assign in_chan_dep_vld_vec_22[23] = dep_chan_vld_27_22;
    assign in_chan_dep_data_vec_22[959 : 920] = dep_chan_data_27_22;
    assign token_in_vec_22[23] = token_27_22;
    assign in_chan_dep_vld_vec_22[24] = dep_chan_vld_28_22;
    assign in_chan_dep_data_vec_22[999 : 960] = dep_chan_data_28_22;
    assign token_in_vec_22[24] = token_28_22;
    assign in_chan_dep_vld_vec_22[25] = dep_chan_vld_29_22;
    assign in_chan_dep_data_vec_22[1039 : 1000] = dep_chan_data_29_22;
    assign token_in_vec_22[25] = token_29_22;
    assign in_chan_dep_vld_vec_22[26] = dep_chan_vld_30_22;
    assign in_chan_dep_data_vec_22[1079 : 1040] = dep_chan_data_30_22;
    assign token_in_vec_22[26] = token_30_22;
    assign in_chan_dep_vld_vec_22[27] = dep_chan_vld_31_22;
    assign in_chan_dep_data_vec_22[1119 : 1080] = dep_chan_data_31_22;
    assign token_in_vec_22[27] = token_31_22;
    assign in_chan_dep_vld_vec_22[28] = dep_chan_vld_32_22;
    assign in_chan_dep_data_vec_22[1159 : 1120] = dep_chan_data_32_22;
    assign token_in_vec_22[28] = token_32_22;
    assign in_chan_dep_vld_vec_22[29] = dep_chan_vld_33_22;
    assign in_chan_dep_data_vec_22[1199 : 1160] = dep_chan_data_33_22;
    assign token_in_vec_22[29] = token_33_22;
    assign in_chan_dep_vld_vec_22[30] = dep_chan_vld_34_22;
    assign in_chan_dep_data_vec_22[1239 : 1200] = dep_chan_data_34_22;
    assign token_in_vec_22[30] = token_34_22;
    assign in_chan_dep_vld_vec_22[31] = dep_chan_vld_35_22;
    assign in_chan_dep_data_vec_22[1279 : 1240] = dep_chan_data_35_22;
    assign token_in_vec_22[31] = token_35_22;
    assign in_chan_dep_vld_vec_22[32] = dep_chan_vld_36_22;
    assign in_chan_dep_data_vec_22[1319 : 1280] = dep_chan_data_36_22;
    assign token_in_vec_22[32] = token_36_22;
    assign dep_chan_vld_22_21 = out_chan_dep_vld_vec_22[0];
    assign dep_chan_data_22_21 = out_chan_dep_data_22;
    assign token_22_21 = token_out_vec_22[0];
    assign dep_chan_vld_22_23 = out_chan_dep_vld_vec_22[1];
    assign dep_chan_data_22_23 = out_chan_dep_data_22;
    assign token_22_23 = token_out_vec_22[1];
    assign dep_chan_vld_22_0 = out_chan_dep_vld_vec_22[2];
    assign dep_chan_data_22_0 = out_chan_dep_data_22;
    assign token_22_0 = token_out_vec_22[2];
    assign dep_chan_vld_22_1 = out_chan_dep_vld_vec_22[3];
    assign dep_chan_data_22_1 = out_chan_dep_data_22;
    assign token_22_1 = token_out_vec_22[3];
    assign dep_chan_vld_22_3 = out_chan_dep_vld_vec_22[4];
    assign dep_chan_data_22_3 = out_chan_dep_data_22;
    assign token_22_3 = token_out_vec_22[4];
    assign dep_chan_vld_22_6 = out_chan_dep_vld_vec_22[5];
    assign dep_chan_data_22_6 = out_chan_dep_data_22;
    assign token_22_6 = token_out_vec_22[5];
    assign dep_chan_vld_22_7 = out_chan_dep_vld_vec_22[6];
    assign dep_chan_data_22_7 = out_chan_dep_data_22;
    assign token_22_7 = token_out_vec_22[6];
    assign dep_chan_vld_22_8 = out_chan_dep_vld_vec_22[7];
    assign dep_chan_data_22_8 = out_chan_dep_data_22;
    assign token_22_8 = token_out_vec_22[7];
    assign dep_chan_vld_22_9 = out_chan_dep_vld_vec_22[8];
    assign dep_chan_data_22_9 = out_chan_dep_data_22;
    assign token_22_9 = token_out_vec_22[8];
    assign dep_chan_vld_22_10 = out_chan_dep_vld_vec_22[9];
    assign dep_chan_data_22_10 = out_chan_dep_data_22;
    assign token_22_10 = token_out_vec_22[9];
    assign dep_chan_vld_22_11 = out_chan_dep_vld_vec_22[10];
    assign dep_chan_data_22_11 = out_chan_dep_data_22;
    assign token_22_11 = token_out_vec_22[10];
    assign dep_chan_vld_22_12 = out_chan_dep_vld_vec_22[11];
    assign dep_chan_data_22_12 = out_chan_dep_data_22;
    assign token_22_12 = token_out_vec_22[11];
    assign dep_chan_vld_22_13 = out_chan_dep_vld_vec_22[12];
    assign dep_chan_data_22_13 = out_chan_dep_data_22;
    assign token_22_13 = token_out_vec_22[12];
    assign dep_chan_vld_22_14 = out_chan_dep_vld_vec_22[13];
    assign dep_chan_data_22_14 = out_chan_dep_data_22;
    assign token_22_14 = token_out_vec_22[13];
    assign dep_chan_vld_22_15 = out_chan_dep_vld_vec_22[14];
    assign dep_chan_data_22_15 = out_chan_dep_data_22;
    assign token_22_15 = token_out_vec_22[14];
    assign dep_chan_vld_22_16 = out_chan_dep_vld_vec_22[15];
    assign dep_chan_data_22_16 = out_chan_dep_data_22;
    assign token_22_16 = token_out_vec_22[15];
    assign dep_chan_vld_22_17 = out_chan_dep_vld_vec_22[16];
    assign dep_chan_data_22_17 = out_chan_dep_data_22;
    assign token_22_17 = token_out_vec_22[16];
    assign dep_chan_vld_22_18 = out_chan_dep_vld_vec_22[17];
    assign dep_chan_data_22_18 = out_chan_dep_data_22;
    assign token_22_18 = token_out_vec_22[17];
    assign dep_chan_vld_22_19 = out_chan_dep_vld_vec_22[18];
    assign dep_chan_data_22_19 = out_chan_dep_data_22;
    assign token_22_19 = token_out_vec_22[18];
    assign dep_chan_vld_22_20 = out_chan_dep_vld_vec_22[19];
    assign dep_chan_data_22_20 = out_chan_dep_data_22;
    assign token_22_20 = token_out_vec_22[19];
    assign dep_chan_vld_22_24 = out_chan_dep_vld_vec_22[20];
    assign dep_chan_data_22_24 = out_chan_dep_data_22;
    assign token_22_24 = token_out_vec_22[20];
    assign dep_chan_vld_22_25 = out_chan_dep_vld_vec_22[21];
    assign dep_chan_data_22_25 = out_chan_dep_data_22;
    assign token_22_25 = token_out_vec_22[21];
    assign dep_chan_vld_22_26 = out_chan_dep_vld_vec_22[22];
    assign dep_chan_data_22_26 = out_chan_dep_data_22;
    assign token_22_26 = token_out_vec_22[22];
    assign dep_chan_vld_22_27 = out_chan_dep_vld_vec_22[23];
    assign dep_chan_data_22_27 = out_chan_dep_data_22;
    assign token_22_27 = token_out_vec_22[23];
    assign dep_chan_vld_22_28 = out_chan_dep_vld_vec_22[24];
    assign dep_chan_data_22_28 = out_chan_dep_data_22;
    assign token_22_28 = token_out_vec_22[24];
    assign dep_chan_vld_22_29 = out_chan_dep_vld_vec_22[25];
    assign dep_chan_data_22_29 = out_chan_dep_data_22;
    assign token_22_29 = token_out_vec_22[25];
    assign dep_chan_vld_22_30 = out_chan_dep_vld_vec_22[26];
    assign dep_chan_data_22_30 = out_chan_dep_data_22;
    assign token_22_30 = token_out_vec_22[26];
    assign dep_chan_vld_22_31 = out_chan_dep_vld_vec_22[27];
    assign dep_chan_data_22_31 = out_chan_dep_data_22;
    assign token_22_31 = token_out_vec_22[27];
    assign dep_chan_vld_22_32 = out_chan_dep_vld_vec_22[28];
    assign dep_chan_data_22_32 = out_chan_dep_data_22;
    assign token_22_32 = token_out_vec_22[28];
    assign dep_chan_vld_22_33 = out_chan_dep_vld_vec_22[29];
    assign dep_chan_data_22_33 = out_chan_dep_data_22;
    assign token_22_33 = token_out_vec_22[29];
    assign dep_chan_vld_22_34 = out_chan_dep_vld_vec_22[30];
    assign dep_chan_data_22_34 = out_chan_dep_data_22;
    assign token_22_34 = token_out_vec_22[30];
    assign dep_chan_vld_22_35 = out_chan_dep_vld_vec_22[31];
    assign dep_chan_data_22_35 = out_chan_dep_data_22;
    assign token_22_35 = token_out_vec_22[31];
    assign dep_chan_vld_22_36 = out_chan_dep_vld_vec_22[32];
    assign dep_chan_data_22_36 = out_chan_dep_data_22;
    assign token_22_36 = token_out_vec_22[32];

    // Process: ProcessingElement_18_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 23, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_23 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_23),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_23),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_23),
        .token_in_vec(token_in_vec_23),
        .dl_detect_in(dl_detect_out),
        .origin(origin[23]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_23),
        .out_chan_dep_data(out_chan_dep_data_23),
        .token_out_vec(token_out_vec_23),
        .dl_detect_out(dl_in_vec[23]));

    assign proc_23_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_17_blk_n) | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_17_blk_n) | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_WriteC_Flattened_fu_179.cPipes_17_blk_n);
    assign proc_23_data_PIPO_blk[0] = 1'b0;
    assign proc_23_start_FIFO_blk[0] = 1'b0;
    assign proc_23_TLF_FIFO_blk[0] = 1'b0;
    assign proc_23_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_23_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_23[0] = dl_detect_out ? proc_dep_vld_vec_23_reg[0] : (proc_23_data_FIFO_blk[0] | proc_23_data_PIPO_blk[0] | proc_23_start_FIFO_blk[0] | proc_23_TLF_FIFO_blk[0] | proc_23_input_sync_blk[0] | proc_23_output_sync_blk[0]);
    assign proc_23_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_18_blk_n) | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_18_blk_n) | (~ProcessingElement_18_U0.grp_ProcessingElement_18_Pipeline_WriteC_Flattened_fu_179.cPipes_18_blk_n);
    assign proc_23_data_PIPO_blk[1] = 1'b0;
    assign proc_23_start_FIFO_blk[1] = 1'b0;
    assign proc_23_TLF_FIFO_blk[1] = 1'b0;
    assign proc_23_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_23_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_23[1] = dl_detect_out ? proc_dep_vld_vec_23_reg[1] : (proc_23_data_FIFO_blk[1] | proc_23_data_PIPO_blk[1] | proc_23_start_FIFO_blk[1] | proc_23_TLF_FIFO_blk[1] | proc_23_input_sync_blk[1] | proc_23_output_sync_blk[1]);
    assign proc_23_data_FIFO_blk[2] = 1'b0;
    assign proc_23_data_PIPO_blk[2] = 1'b0;
    assign proc_23_start_FIFO_blk[2] = 1'b0;
    assign proc_23_TLF_FIFO_blk[2] = 1'b0;
    assign proc_23_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_23_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_23[2] = dl_detect_out ? proc_dep_vld_vec_23_reg[2] : (proc_23_data_FIFO_blk[2] | proc_23_data_PIPO_blk[2] | proc_23_start_FIFO_blk[2] | proc_23_TLF_FIFO_blk[2] | proc_23_input_sync_blk[2] | proc_23_output_sync_blk[2]);
    assign proc_23_data_FIFO_blk[3] = 1'b0;
    assign proc_23_data_PIPO_blk[3] = 1'b0;
    assign proc_23_start_FIFO_blk[3] = 1'b0;
    assign proc_23_TLF_FIFO_blk[3] = 1'b0;
    assign proc_23_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_23_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_23[3] = dl_detect_out ? proc_dep_vld_vec_23_reg[3] : (proc_23_data_FIFO_blk[3] | proc_23_data_PIPO_blk[3] | proc_23_start_FIFO_blk[3] | proc_23_TLF_FIFO_blk[3] | proc_23_input_sync_blk[3] | proc_23_output_sync_blk[3]);
    assign proc_23_data_FIFO_blk[4] = 1'b0;
    assign proc_23_data_PIPO_blk[4] = 1'b0;
    assign proc_23_start_FIFO_blk[4] = 1'b0;
    assign proc_23_TLF_FIFO_blk[4] = 1'b0;
    assign proc_23_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_23_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_23[4] = dl_detect_out ? proc_dep_vld_vec_23_reg[4] : (proc_23_data_FIFO_blk[4] | proc_23_data_PIPO_blk[4] | proc_23_start_FIFO_blk[4] | proc_23_TLF_FIFO_blk[4] | proc_23_input_sync_blk[4] | proc_23_output_sync_blk[4]);
    assign proc_23_data_FIFO_blk[5] = 1'b0;
    assign proc_23_data_PIPO_blk[5] = 1'b0;
    assign proc_23_start_FIFO_blk[5] = 1'b0;
    assign proc_23_TLF_FIFO_blk[5] = 1'b0;
    assign proc_23_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_23_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_23[5] = dl_detect_out ? proc_dep_vld_vec_23_reg[5] : (proc_23_data_FIFO_blk[5] | proc_23_data_PIPO_blk[5] | proc_23_start_FIFO_blk[5] | proc_23_TLF_FIFO_blk[5] | proc_23_input_sync_blk[5] | proc_23_output_sync_blk[5]);
    assign proc_23_data_FIFO_blk[6] = 1'b0;
    assign proc_23_data_PIPO_blk[6] = 1'b0;
    assign proc_23_start_FIFO_blk[6] = 1'b0;
    assign proc_23_TLF_FIFO_blk[6] = 1'b0;
    assign proc_23_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_23_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_23[6] = dl_detect_out ? proc_dep_vld_vec_23_reg[6] : (proc_23_data_FIFO_blk[6] | proc_23_data_PIPO_blk[6] | proc_23_start_FIFO_blk[6] | proc_23_TLF_FIFO_blk[6] | proc_23_input_sync_blk[6] | proc_23_output_sync_blk[6]);
    assign proc_23_data_FIFO_blk[7] = 1'b0;
    assign proc_23_data_PIPO_blk[7] = 1'b0;
    assign proc_23_start_FIFO_blk[7] = 1'b0;
    assign proc_23_TLF_FIFO_blk[7] = 1'b0;
    assign proc_23_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_23_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_23[7] = dl_detect_out ? proc_dep_vld_vec_23_reg[7] : (proc_23_data_FIFO_blk[7] | proc_23_data_PIPO_blk[7] | proc_23_start_FIFO_blk[7] | proc_23_TLF_FIFO_blk[7] | proc_23_input_sync_blk[7] | proc_23_output_sync_blk[7]);
    assign proc_23_data_FIFO_blk[8] = 1'b0;
    assign proc_23_data_PIPO_blk[8] = 1'b0;
    assign proc_23_start_FIFO_blk[8] = 1'b0;
    assign proc_23_TLF_FIFO_blk[8] = 1'b0;
    assign proc_23_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_23_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_23[8] = dl_detect_out ? proc_dep_vld_vec_23_reg[8] : (proc_23_data_FIFO_blk[8] | proc_23_data_PIPO_blk[8] | proc_23_start_FIFO_blk[8] | proc_23_TLF_FIFO_blk[8] | proc_23_input_sync_blk[8] | proc_23_output_sync_blk[8]);
    assign proc_23_data_FIFO_blk[9] = 1'b0;
    assign proc_23_data_PIPO_blk[9] = 1'b0;
    assign proc_23_start_FIFO_blk[9] = 1'b0;
    assign proc_23_TLF_FIFO_blk[9] = 1'b0;
    assign proc_23_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_23_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_23[9] = dl_detect_out ? proc_dep_vld_vec_23_reg[9] : (proc_23_data_FIFO_blk[9] | proc_23_data_PIPO_blk[9] | proc_23_start_FIFO_blk[9] | proc_23_TLF_FIFO_blk[9] | proc_23_input_sync_blk[9] | proc_23_output_sync_blk[9]);
    assign proc_23_data_FIFO_blk[10] = 1'b0;
    assign proc_23_data_PIPO_blk[10] = 1'b0;
    assign proc_23_start_FIFO_blk[10] = 1'b0;
    assign proc_23_TLF_FIFO_blk[10] = 1'b0;
    assign proc_23_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_23_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_23[10] = dl_detect_out ? proc_dep_vld_vec_23_reg[10] : (proc_23_data_FIFO_blk[10] | proc_23_data_PIPO_blk[10] | proc_23_start_FIFO_blk[10] | proc_23_TLF_FIFO_blk[10] | proc_23_input_sync_blk[10] | proc_23_output_sync_blk[10]);
    assign proc_23_data_FIFO_blk[11] = 1'b0;
    assign proc_23_data_PIPO_blk[11] = 1'b0;
    assign proc_23_start_FIFO_blk[11] = 1'b0;
    assign proc_23_TLF_FIFO_blk[11] = 1'b0;
    assign proc_23_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_23_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_23[11] = dl_detect_out ? proc_dep_vld_vec_23_reg[11] : (proc_23_data_FIFO_blk[11] | proc_23_data_PIPO_blk[11] | proc_23_start_FIFO_blk[11] | proc_23_TLF_FIFO_blk[11] | proc_23_input_sync_blk[11] | proc_23_output_sync_blk[11]);
    assign proc_23_data_FIFO_blk[12] = 1'b0;
    assign proc_23_data_PIPO_blk[12] = 1'b0;
    assign proc_23_start_FIFO_blk[12] = 1'b0;
    assign proc_23_TLF_FIFO_blk[12] = 1'b0;
    assign proc_23_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_23_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_23[12] = dl_detect_out ? proc_dep_vld_vec_23_reg[12] : (proc_23_data_FIFO_blk[12] | proc_23_data_PIPO_blk[12] | proc_23_start_FIFO_blk[12] | proc_23_TLF_FIFO_blk[12] | proc_23_input_sync_blk[12] | proc_23_output_sync_blk[12]);
    assign proc_23_data_FIFO_blk[13] = 1'b0;
    assign proc_23_data_PIPO_blk[13] = 1'b0;
    assign proc_23_start_FIFO_blk[13] = 1'b0;
    assign proc_23_TLF_FIFO_blk[13] = 1'b0;
    assign proc_23_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_23_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_23[13] = dl_detect_out ? proc_dep_vld_vec_23_reg[13] : (proc_23_data_FIFO_blk[13] | proc_23_data_PIPO_blk[13] | proc_23_start_FIFO_blk[13] | proc_23_TLF_FIFO_blk[13] | proc_23_input_sync_blk[13] | proc_23_output_sync_blk[13]);
    assign proc_23_data_FIFO_blk[14] = 1'b0;
    assign proc_23_data_PIPO_blk[14] = 1'b0;
    assign proc_23_start_FIFO_blk[14] = 1'b0;
    assign proc_23_TLF_FIFO_blk[14] = 1'b0;
    assign proc_23_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_23_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_23[14] = dl_detect_out ? proc_dep_vld_vec_23_reg[14] : (proc_23_data_FIFO_blk[14] | proc_23_data_PIPO_blk[14] | proc_23_start_FIFO_blk[14] | proc_23_TLF_FIFO_blk[14] | proc_23_input_sync_blk[14] | proc_23_output_sync_blk[14]);
    assign proc_23_data_FIFO_blk[15] = 1'b0;
    assign proc_23_data_PIPO_blk[15] = 1'b0;
    assign proc_23_start_FIFO_blk[15] = 1'b0;
    assign proc_23_TLF_FIFO_blk[15] = 1'b0;
    assign proc_23_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_23_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_23[15] = dl_detect_out ? proc_dep_vld_vec_23_reg[15] : (proc_23_data_FIFO_blk[15] | proc_23_data_PIPO_blk[15] | proc_23_start_FIFO_blk[15] | proc_23_TLF_FIFO_blk[15] | proc_23_input_sync_blk[15] | proc_23_output_sync_blk[15]);
    assign proc_23_data_FIFO_blk[16] = 1'b0;
    assign proc_23_data_PIPO_blk[16] = 1'b0;
    assign proc_23_start_FIFO_blk[16] = 1'b0;
    assign proc_23_TLF_FIFO_blk[16] = 1'b0;
    assign proc_23_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_23_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_23[16] = dl_detect_out ? proc_dep_vld_vec_23_reg[16] : (proc_23_data_FIFO_blk[16] | proc_23_data_PIPO_blk[16] | proc_23_start_FIFO_blk[16] | proc_23_TLF_FIFO_blk[16] | proc_23_input_sync_blk[16] | proc_23_output_sync_blk[16]);
    assign proc_23_data_FIFO_blk[17] = 1'b0;
    assign proc_23_data_PIPO_blk[17] = 1'b0;
    assign proc_23_start_FIFO_blk[17] = 1'b0;
    assign proc_23_TLF_FIFO_blk[17] = 1'b0;
    assign proc_23_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_23_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_23[17] = dl_detect_out ? proc_dep_vld_vec_23_reg[17] : (proc_23_data_FIFO_blk[17] | proc_23_data_PIPO_blk[17] | proc_23_start_FIFO_blk[17] | proc_23_TLF_FIFO_blk[17] | proc_23_input_sync_blk[17] | proc_23_output_sync_blk[17]);
    assign proc_23_data_FIFO_blk[18] = 1'b0;
    assign proc_23_data_PIPO_blk[18] = 1'b0;
    assign proc_23_start_FIFO_blk[18] = 1'b0;
    assign proc_23_TLF_FIFO_blk[18] = 1'b0;
    assign proc_23_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_23_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_23[18] = dl_detect_out ? proc_dep_vld_vec_23_reg[18] : (proc_23_data_FIFO_blk[18] | proc_23_data_PIPO_blk[18] | proc_23_start_FIFO_blk[18] | proc_23_TLF_FIFO_blk[18] | proc_23_input_sync_blk[18] | proc_23_output_sync_blk[18]);
    assign proc_23_data_FIFO_blk[19] = 1'b0;
    assign proc_23_data_PIPO_blk[19] = 1'b0;
    assign proc_23_start_FIFO_blk[19] = 1'b0;
    assign proc_23_TLF_FIFO_blk[19] = 1'b0;
    assign proc_23_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_23_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_23[19] = dl_detect_out ? proc_dep_vld_vec_23_reg[19] : (proc_23_data_FIFO_blk[19] | proc_23_data_PIPO_blk[19] | proc_23_start_FIFO_blk[19] | proc_23_TLF_FIFO_blk[19] | proc_23_input_sync_blk[19] | proc_23_output_sync_blk[19]);
    assign proc_23_data_FIFO_blk[20] = 1'b0;
    assign proc_23_data_PIPO_blk[20] = 1'b0;
    assign proc_23_start_FIFO_blk[20] = 1'b0;
    assign proc_23_TLF_FIFO_blk[20] = 1'b0;
    assign proc_23_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_23_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_23[20] = dl_detect_out ? proc_dep_vld_vec_23_reg[20] : (proc_23_data_FIFO_blk[20] | proc_23_data_PIPO_blk[20] | proc_23_start_FIFO_blk[20] | proc_23_TLF_FIFO_blk[20] | proc_23_input_sync_blk[20] | proc_23_output_sync_blk[20]);
    assign proc_23_data_FIFO_blk[21] = 1'b0;
    assign proc_23_data_PIPO_blk[21] = 1'b0;
    assign proc_23_start_FIFO_blk[21] = 1'b0;
    assign proc_23_TLF_FIFO_blk[21] = 1'b0;
    assign proc_23_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_23_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_23[21] = dl_detect_out ? proc_dep_vld_vec_23_reg[21] : (proc_23_data_FIFO_blk[21] | proc_23_data_PIPO_blk[21] | proc_23_start_FIFO_blk[21] | proc_23_TLF_FIFO_blk[21] | proc_23_input_sync_blk[21] | proc_23_output_sync_blk[21]);
    assign proc_23_data_FIFO_blk[22] = 1'b0;
    assign proc_23_data_PIPO_blk[22] = 1'b0;
    assign proc_23_start_FIFO_blk[22] = 1'b0;
    assign proc_23_TLF_FIFO_blk[22] = 1'b0;
    assign proc_23_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_23_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_23[22] = dl_detect_out ? proc_dep_vld_vec_23_reg[22] : (proc_23_data_FIFO_blk[22] | proc_23_data_PIPO_blk[22] | proc_23_start_FIFO_blk[22] | proc_23_TLF_FIFO_blk[22] | proc_23_input_sync_blk[22] | proc_23_output_sync_blk[22]);
    assign proc_23_data_FIFO_blk[23] = 1'b0;
    assign proc_23_data_PIPO_blk[23] = 1'b0;
    assign proc_23_start_FIFO_blk[23] = 1'b0;
    assign proc_23_TLF_FIFO_blk[23] = 1'b0;
    assign proc_23_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_23_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_23[23] = dl_detect_out ? proc_dep_vld_vec_23_reg[23] : (proc_23_data_FIFO_blk[23] | proc_23_data_PIPO_blk[23] | proc_23_start_FIFO_blk[23] | proc_23_TLF_FIFO_blk[23] | proc_23_input_sync_blk[23] | proc_23_output_sync_blk[23]);
    assign proc_23_data_FIFO_blk[24] = 1'b0;
    assign proc_23_data_PIPO_blk[24] = 1'b0;
    assign proc_23_start_FIFO_blk[24] = 1'b0;
    assign proc_23_TLF_FIFO_blk[24] = 1'b0;
    assign proc_23_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_23_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_23[24] = dl_detect_out ? proc_dep_vld_vec_23_reg[24] : (proc_23_data_FIFO_blk[24] | proc_23_data_PIPO_blk[24] | proc_23_start_FIFO_blk[24] | proc_23_TLF_FIFO_blk[24] | proc_23_input_sync_blk[24] | proc_23_output_sync_blk[24]);
    assign proc_23_data_FIFO_blk[25] = 1'b0;
    assign proc_23_data_PIPO_blk[25] = 1'b0;
    assign proc_23_start_FIFO_blk[25] = 1'b0;
    assign proc_23_TLF_FIFO_blk[25] = 1'b0;
    assign proc_23_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_23_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_23[25] = dl_detect_out ? proc_dep_vld_vec_23_reg[25] : (proc_23_data_FIFO_blk[25] | proc_23_data_PIPO_blk[25] | proc_23_start_FIFO_blk[25] | proc_23_TLF_FIFO_blk[25] | proc_23_input_sync_blk[25] | proc_23_output_sync_blk[25]);
    assign proc_23_data_FIFO_blk[26] = 1'b0;
    assign proc_23_data_PIPO_blk[26] = 1'b0;
    assign proc_23_start_FIFO_blk[26] = 1'b0;
    assign proc_23_TLF_FIFO_blk[26] = 1'b0;
    assign proc_23_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_23_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_23[26] = dl_detect_out ? proc_dep_vld_vec_23_reg[26] : (proc_23_data_FIFO_blk[26] | proc_23_data_PIPO_blk[26] | proc_23_start_FIFO_blk[26] | proc_23_TLF_FIFO_blk[26] | proc_23_input_sync_blk[26] | proc_23_output_sync_blk[26]);
    assign proc_23_data_FIFO_blk[27] = 1'b0;
    assign proc_23_data_PIPO_blk[27] = 1'b0;
    assign proc_23_start_FIFO_blk[27] = 1'b0;
    assign proc_23_TLF_FIFO_blk[27] = 1'b0;
    assign proc_23_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_23_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_23[27] = dl_detect_out ? proc_dep_vld_vec_23_reg[27] : (proc_23_data_FIFO_blk[27] | proc_23_data_PIPO_blk[27] | proc_23_start_FIFO_blk[27] | proc_23_TLF_FIFO_blk[27] | proc_23_input_sync_blk[27] | proc_23_output_sync_blk[27]);
    assign proc_23_data_FIFO_blk[28] = 1'b0;
    assign proc_23_data_PIPO_blk[28] = 1'b0;
    assign proc_23_start_FIFO_blk[28] = 1'b0;
    assign proc_23_TLF_FIFO_blk[28] = 1'b0;
    assign proc_23_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_23_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_23[28] = dl_detect_out ? proc_dep_vld_vec_23_reg[28] : (proc_23_data_FIFO_blk[28] | proc_23_data_PIPO_blk[28] | proc_23_start_FIFO_blk[28] | proc_23_TLF_FIFO_blk[28] | proc_23_input_sync_blk[28] | proc_23_output_sync_blk[28]);
    assign proc_23_data_FIFO_blk[29] = 1'b0;
    assign proc_23_data_PIPO_blk[29] = 1'b0;
    assign proc_23_start_FIFO_blk[29] = 1'b0;
    assign proc_23_TLF_FIFO_blk[29] = 1'b0;
    assign proc_23_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_23_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_23[29] = dl_detect_out ? proc_dep_vld_vec_23_reg[29] : (proc_23_data_FIFO_blk[29] | proc_23_data_PIPO_blk[29] | proc_23_start_FIFO_blk[29] | proc_23_TLF_FIFO_blk[29] | proc_23_input_sync_blk[29] | proc_23_output_sync_blk[29]);
    assign proc_23_data_FIFO_blk[30] = 1'b0;
    assign proc_23_data_PIPO_blk[30] = 1'b0;
    assign proc_23_start_FIFO_blk[30] = 1'b0;
    assign proc_23_TLF_FIFO_blk[30] = 1'b0;
    assign proc_23_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_23_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_23[30] = dl_detect_out ? proc_dep_vld_vec_23_reg[30] : (proc_23_data_FIFO_blk[30] | proc_23_data_PIPO_blk[30] | proc_23_start_FIFO_blk[30] | proc_23_TLF_FIFO_blk[30] | proc_23_input_sync_blk[30] | proc_23_output_sync_blk[30]);
    assign proc_23_data_FIFO_blk[31] = 1'b0;
    assign proc_23_data_PIPO_blk[31] = 1'b0;
    assign proc_23_start_FIFO_blk[31] = 1'b0;
    assign proc_23_TLF_FIFO_blk[31] = 1'b0;
    assign proc_23_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_23_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_23[31] = dl_detect_out ? proc_dep_vld_vec_23_reg[31] : (proc_23_data_FIFO_blk[31] | proc_23_data_PIPO_blk[31] | proc_23_start_FIFO_blk[31] | proc_23_TLF_FIFO_blk[31] | proc_23_input_sync_blk[31] | proc_23_output_sync_blk[31]);
    assign proc_23_data_FIFO_blk[32] = 1'b0;
    assign proc_23_data_PIPO_blk[32] = 1'b0;
    assign proc_23_start_FIFO_blk[32] = 1'b0;
    assign proc_23_TLF_FIFO_blk[32] = 1'b0;
    assign proc_23_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_18_U0_ap_ready & ProcessingElement_18_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_23_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_23[32] = dl_detect_out ? proc_dep_vld_vec_23_reg[32] : (proc_23_data_FIFO_blk[32] | proc_23_data_PIPO_blk[32] | proc_23_start_FIFO_blk[32] | proc_23_TLF_FIFO_blk[32] | proc_23_input_sync_blk[32] | proc_23_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_23_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_23_reg <= proc_dep_vld_vec_23;
        end
    end
    assign in_chan_dep_vld_vec_23[0] = dep_chan_vld_0_23;
    assign in_chan_dep_data_vec_23[39 : 0] = dep_chan_data_0_23;
    assign token_in_vec_23[0] = token_0_23;
    assign in_chan_dep_vld_vec_23[1] = dep_chan_vld_1_23;
    assign in_chan_dep_data_vec_23[79 : 40] = dep_chan_data_1_23;
    assign token_in_vec_23[1] = token_1_23;
    assign in_chan_dep_vld_vec_23[2] = dep_chan_vld_3_23;
    assign in_chan_dep_data_vec_23[119 : 80] = dep_chan_data_3_23;
    assign token_in_vec_23[2] = token_3_23;
    assign in_chan_dep_vld_vec_23[3] = dep_chan_vld_6_23;
    assign in_chan_dep_data_vec_23[159 : 120] = dep_chan_data_6_23;
    assign token_in_vec_23[3] = token_6_23;
    assign in_chan_dep_vld_vec_23[4] = dep_chan_vld_7_23;
    assign in_chan_dep_data_vec_23[199 : 160] = dep_chan_data_7_23;
    assign token_in_vec_23[4] = token_7_23;
    assign in_chan_dep_vld_vec_23[5] = dep_chan_vld_8_23;
    assign in_chan_dep_data_vec_23[239 : 200] = dep_chan_data_8_23;
    assign token_in_vec_23[5] = token_8_23;
    assign in_chan_dep_vld_vec_23[6] = dep_chan_vld_9_23;
    assign in_chan_dep_data_vec_23[279 : 240] = dep_chan_data_9_23;
    assign token_in_vec_23[6] = token_9_23;
    assign in_chan_dep_vld_vec_23[7] = dep_chan_vld_10_23;
    assign in_chan_dep_data_vec_23[319 : 280] = dep_chan_data_10_23;
    assign token_in_vec_23[7] = token_10_23;
    assign in_chan_dep_vld_vec_23[8] = dep_chan_vld_11_23;
    assign in_chan_dep_data_vec_23[359 : 320] = dep_chan_data_11_23;
    assign token_in_vec_23[8] = token_11_23;
    assign in_chan_dep_vld_vec_23[9] = dep_chan_vld_12_23;
    assign in_chan_dep_data_vec_23[399 : 360] = dep_chan_data_12_23;
    assign token_in_vec_23[9] = token_12_23;
    assign in_chan_dep_vld_vec_23[10] = dep_chan_vld_13_23;
    assign in_chan_dep_data_vec_23[439 : 400] = dep_chan_data_13_23;
    assign token_in_vec_23[10] = token_13_23;
    assign in_chan_dep_vld_vec_23[11] = dep_chan_vld_14_23;
    assign in_chan_dep_data_vec_23[479 : 440] = dep_chan_data_14_23;
    assign token_in_vec_23[11] = token_14_23;
    assign in_chan_dep_vld_vec_23[12] = dep_chan_vld_15_23;
    assign in_chan_dep_data_vec_23[519 : 480] = dep_chan_data_15_23;
    assign token_in_vec_23[12] = token_15_23;
    assign in_chan_dep_vld_vec_23[13] = dep_chan_vld_16_23;
    assign in_chan_dep_data_vec_23[559 : 520] = dep_chan_data_16_23;
    assign token_in_vec_23[13] = token_16_23;
    assign in_chan_dep_vld_vec_23[14] = dep_chan_vld_17_23;
    assign in_chan_dep_data_vec_23[599 : 560] = dep_chan_data_17_23;
    assign token_in_vec_23[14] = token_17_23;
    assign in_chan_dep_vld_vec_23[15] = dep_chan_vld_18_23;
    assign in_chan_dep_data_vec_23[639 : 600] = dep_chan_data_18_23;
    assign token_in_vec_23[15] = token_18_23;
    assign in_chan_dep_vld_vec_23[16] = dep_chan_vld_19_23;
    assign in_chan_dep_data_vec_23[679 : 640] = dep_chan_data_19_23;
    assign token_in_vec_23[16] = token_19_23;
    assign in_chan_dep_vld_vec_23[17] = dep_chan_vld_20_23;
    assign in_chan_dep_data_vec_23[719 : 680] = dep_chan_data_20_23;
    assign token_in_vec_23[17] = token_20_23;
    assign in_chan_dep_vld_vec_23[18] = dep_chan_vld_21_23;
    assign in_chan_dep_data_vec_23[759 : 720] = dep_chan_data_21_23;
    assign token_in_vec_23[18] = token_21_23;
    assign in_chan_dep_vld_vec_23[19] = dep_chan_vld_22_23;
    assign in_chan_dep_data_vec_23[799 : 760] = dep_chan_data_22_23;
    assign token_in_vec_23[19] = token_22_23;
    assign in_chan_dep_vld_vec_23[20] = dep_chan_vld_24_23;
    assign in_chan_dep_data_vec_23[839 : 800] = dep_chan_data_24_23;
    assign token_in_vec_23[20] = token_24_23;
    assign in_chan_dep_vld_vec_23[21] = dep_chan_vld_25_23;
    assign in_chan_dep_data_vec_23[879 : 840] = dep_chan_data_25_23;
    assign token_in_vec_23[21] = token_25_23;
    assign in_chan_dep_vld_vec_23[22] = dep_chan_vld_26_23;
    assign in_chan_dep_data_vec_23[919 : 880] = dep_chan_data_26_23;
    assign token_in_vec_23[22] = token_26_23;
    assign in_chan_dep_vld_vec_23[23] = dep_chan_vld_27_23;
    assign in_chan_dep_data_vec_23[959 : 920] = dep_chan_data_27_23;
    assign token_in_vec_23[23] = token_27_23;
    assign in_chan_dep_vld_vec_23[24] = dep_chan_vld_28_23;
    assign in_chan_dep_data_vec_23[999 : 960] = dep_chan_data_28_23;
    assign token_in_vec_23[24] = token_28_23;
    assign in_chan_dep_vld_vec_23[25] = dep_chan_vld_29_23;
    assign in_chan_dep_data_vec_23[1039 : 1000] = dep_chan_data_29_23;
    assign token_in_vec_23[25] = token_29_23;
    assign in_chan_dep_vld_vec_23[26] = dep_chan_vld_30_23;
    assign in_chan_dep_data_vec_23[1079 : 1040] = dep_chan_data_30_23;
    assign token_in_vec_23[26] = token_30_23;
    assign in_chan_dep_vld_vec_23[27] = dep_chan_vld_31_23;
    assign in_chan_dep_data_vec_23[1119 : 1080] = dep_chan_data_31_23;
    assign token_in_vec_23[27] = token_31_23;
    assign in_chan_dep_vld_vec_23[28] = dep_chan_vld_32_23;
    assign in_chan_dep_data_vec_23[1159 : 1120] = dep_chan_data_32_23;
    assign token_in_vec_23[28] = token_32_23;
    assign in_chan_dep_vld_vec_23[29] = dep_chan_vld_33_23;
    assign in_chan_dep_data_vec_23[1199 : 1160] = dep_chan_data_33_23;
    assign token_in_vec_23[29] = token_33_23;
    assign in_chan_dep_vld_vec_23[30] = dep_chan_vld_34_23;
    assign in_chan_dep_data_vec_23[1239 : 1200] = dep_chan_data_34_23;
    assign token_in_vec_23[30] = token_34_23;
    assign in_chan_dep_vld_vec_23[31] = dep_chan_vld_35_23;
    assign in_chan_dep_data_vec_23[1279 : 1240] = dep_chan_data_35_23;
    assign token_in_vec_23[31] = token_35_23;
    assign in_chan_dep_vld_vec_23[32] = dep_chan_vld_36_23;
    assign in_chan_dep_data_vec_23[1319 : 1280] = dep_chan_data_36_23;
    assign token_in_vec_23[32] = token_36_23;
    assign dep_chan_vld_23_22 = out_chan_dep_vld_vec_23[0];
    assign dep_chan_data_23_22 = out_chan_dep_data_23;
    assign token_23_22 = token_out_vec_23[0];
    assign dep_chan_vld_23_24 = out_chan_dep_vld_vec_23[1];
    assign dep_chan_data_23_24 = out_chan_dep_data_23;
    assign token_23_24 = token_out_vec_23[1];
    assign dep_chan_vld_23_0 = out_chan_dep_vld_vec_23[2];
    assign dep_chan_data_23_0 = out_chan_dep_data_23;
    assign token_23_0 = token_out_vec_23[2];
    assign dep_chan_vld_23_1 = out_chan_dep_vld_vec_23[3];
    assign dep_chan_data_23_1 = out_chan_dep_data_23;
    assign token_23_1 = token_out_vec_23[3];
    assign dep_chan_vld_23_3 = out_chan_dep_vld_vec_23[4];
    assign dep_chan_data_23_3 = out_chan_dep_data_23;
    assign token_23_3 = token_out_vec_23[4];
    assign dep_chan_vld_23_6 = out_chan_dep_vld_vec_23[5];
    assign dep_chan_data_23_6 = out_chan_dep_data_23;
    assign token_23_6 = token_out_vec_23[5];
    assign dep_chan_vld_23_7 = out_chan_dep_vld_vec_23[6];
    assign dep_chan_data_23_7 = out_chan_dep_data_23;
    assign token_23_7 = token_out_vec_23[6];
    assign dep_chan_vld_23_8 = out_chan_dep_vld_vec_23[7];
    assign dep_chan_data_23_8 = out_chan_dep_data_23;
    assign token_23_8 = token_out_vec_23[7];
    assign dep_chan_vld_23_9 = out_chan_dep_vld_vec_23[8];
    assign dep_chan_data_23_9 = out_chan_dep_data_23;
    assign token_23_9 = token_out_vec_23[8];
    assign dep_chan_vld_23_10 = out_chan_dep_vld_vec_23[9];
    assign dep_chan_data_23_10 = out_chan_dep_data_23;
    assign token_23_10 = token_out_vec_23[9];
    assign dep_chan_vld_23_11 = out_chan_dep_vld_vec_23[10];
    assign dep_chan_data_23_11 = out_chan_dep_data_23;
    assign token_23_11 = token_out_vec_23[10];
    assign dep_chan_vld_23_12 = out_chan_dep_vld_vec_23[11];
    assign dep_chan_data_23_12 = out_chan_dep_data_23;
    assign token_23_12 = token_out_vec_23[11];
    assign dep_chan_vld_23_13 = out_chan_dep_vld_vec_23[12];
    assign dep_chan_data_23_13 = out_chan_dep_data_23;
    assign token_23_13 = token_out_vec_23[12];
    assign dep_chan_vld_23_14 = out_chan_dep_vld_vec_23[13];
    assign dep_chan_data_23_14 = out_chan_dep_data_23;
    assign token_23_14 = token_out_vec_23[13];
    assign dep_chan_vld_23_15 = out_chan_dep_vld_vec_23[14];
    assign dep_chan_data_23_15 = out_chan_dep_data_23;
    assign token_23_15 = token_out_vec_23[14];
    assign dep_chan_vld_23_16 = out_chan_dep_vld_vec_23[15];
    assign dep_chan_data_23_16 = out_chan_dep_data_23;
    assign token_23_16 = token_out_vec_23[15];
    assign dep_chan_vld_23_17 = out_chan_dep_vld_vec_23[16];
    assign dep_chan_data_23_17 = out_chan_dep_data_23;
    assign token_23_17 = token_out_vec_23[16];
    assign dep_chan_vld_23_18 = out_chan_dep_vld_vec_23[17];
    assign dep_chan_data_23_18 = out_chan_dep_data_23;
    assign token_23_18 = token_out_vec_23[17];
    assign dep_chan_vld_23_19 = out_chan_dep_vld_vec_23[18];
    assign dep_chan_data_23_19 = out_chan_dep_data_23;
    assign token_23_19 = token_out_vec_23[18];
    assign dep_chan_vld_23_20 = out_chan_dep_vld_vec_23[19];
    assign dep_chan_data_23_20 = out_chan_dep_data_23;
    assign token_23_20 = token_out_vec_23[19];
    assign dep_chan_vld_23_21 = out_chan_dep_vld_vec_23[20];
    assign dep_chan_data_23_21 = out_chan_dep_data_23;
    assign token_23_21 = token_out_vec_23[20];
    assign dep_chan_vld_23_25 = out_chan_dep_vld_vec_23[21];
    assign dep_chan_data_23_25 = out_chan_dep_data_23;
    assign token_23_25 = token_out_vec_23[21];
    assign dep_chan_vld_23_26 = out_chan_dep_vld_vec_23[22];
    assign dep_chan_data_23_26 = out_chan_dep_data_23;
    assign token_23_26 = token_out_vec_23[22];
    assign dep_chan_vld_23_27 = out_chan_dep_vld_vec_23[23];
    assign dep_chan_data_23_27 = out_chan_dep_data_23;
    assign token_23_27 = token_out_vec_23[23];
    assign dep_chan_vld_23_28 = out_chan_dep_vld_vec_23[24];
    assign dep_chan_data_23_28 = out_chan_dep_data_23;
    assign token_23_28 = token_out_vec_23[24];
    assign dep_chan_vld_23_29 = out_chan_dep_vld_vec_23[25];
    assign dep_chan_data_23_29 = out_chan_dep_data_23;
    assign token_23_29 = token_out_vec_23[25];
    assign dep_chan_vld_23_30 = out_chan_dep_vld_vec_23[26];
    assign dep_chan_data_23_30 = out_chan_dep_data_23;
    assign token_23_30 = token_out_vec_23[26];
    assign dep_chan_vld_23_31 = out_chan_dep_vld_vec_23[27];
    assign dep_chan_data_23_31 = out_chan_dep_data_23;
    assign token_23_31 = token_out_vec_23[27];
    assign dep_chan_vld_23_32 = out_chan_dep_vld_vec_23[28];
    assign dep_chan_data_23_32 = out_chan_dep_data_23;
    assign token_23_32 = token_out_vec_23[28];
    assign dep_chan_vld_23_33 = out_chan_dep_vld_vec_23[29];
    assign dep_chan_data_23_33 = out_chan_dep_data_23;
    assign token_23_33 = token_out_vec_23[29];
    assign dep_chan_vld_23_34 = out_chan_dep_vld_vec_23[30];
    assign dep_chan_data_23_34 = out_chan_dep_data_23;
    assign token_23_34 = token_out_vec_23[30];
    assign dep_chan_vld_23_35 = out_chan_dep_vld_vec_23[31];
    assign dep_chan_data_23_35 = out_chan_dep_data_23;
    assign token_23_35 = token_out_vec_23[31];
    assign dep_chan_vld_23_36 = out_chan_dep_vld_vec_23[32];
    assign dep_chan_data_23_36 = out_chan_dep_data_23;
    assign token_23_36 = token_out_vec_23[32];

    // Process: ProcessingElement_19_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 24, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_24 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_24),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_24),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_24),
        .token_in_vec(token_in_vec_24),
        .dl_detect_in(dl_detect_out),
        .origin(origin[24]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_24),
        .out_chan_dep_data(out_chan_dep_data_24),
        .token_out_vec(token_out_vec_24),
        .dl_detect_out(dl_in_vec[24]));

    assign proc_24_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_18_blk_n) | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_18_blk_n) | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_WriteC_Flattened_fu_179.cPipes_18_blk_n);
    assign proc_24_data_PIPO_blk[0] = 1'b0;
    assign proc_24_start_FIFO_blk[0] = 1'b0;
    assign proc_24_TLF_FIFO_blk[0] = 1'b0;
    assign proc_24_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_24_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_24[0] = dl_detect_out ? proc_dep_vld_vec_24_reg[0] : (proc_24_data_FIFO_blk[0] | proc_24_data_PIPO_blk[0] | proc_24_start_FIFO_blk[0] | proc_24_TLF_FIFO_blk[0] | proc_24_input_sync_blk[0] | proc_24_output_sync_blk[0]);
    assign proc_24_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_19_blk_n) | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_19_blk_n) | (~ProcessingElement_19_U0.grp_ProcessingElement_19_Pipeline_WriteC_Flattened_fu_179.cPipes_19_blk_n);
    assign proc_24_data_PIPO_blk[1] = 1'b0;
    assign proc_24_start_FIFO_blk[1] = 1'b0;
    assign proc_24_TLF_FIFO_blk[1] = 1'b0;
    assign proc_24_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_24_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_24[1] = dl_detect_out ? proc_dep_vld_vec_24_reg[1] : (proc_24_data_FIFO_blk[1] | proc_24_data_PIPO_blk[1] | proc_24_start_FIFO_blk[1] | proc_24_TLF_FIFO_blk[1] | proc_24_input_sync_blk[1] | proc_24_output_sync_blk[1]);
    assign proc_24_data_FIFO_blk[2] = 1'b0;
    assign proc_24_data_PIPO_blk[2] = 1'b0;
    assign proc_24_start_FIFO_blk[2] = 1'b0;
    assign proc_24_TLF_FIFO_blk[2] = 1'b0;
    assign proc_24_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_24_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_24[2] = dl_detect_out ? proc_dep_vld_vec_24_reg[2] : (proc_24_data_FIFO_blk[2] | proc_24_data_PIPO_blk[2] | proc_24_start_FIFO_blk[2] | proc_24_TLF_FIFO_blk[2] | proc_24_input_sync_blk[2] | proc_24_output_sync_blk[2]);
    assign proc_24_data_FIFO_blk[3] = 1'b0;
    assign proc_24_data_PIPO_blk[3] = 1'b0;
    assign proc_24_start_FIFO_blk[3] = 1'b0;
    assign proc_24_TLF_FIFO_blk[3] = 1'b0;
    assign proc_24_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_24_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_24[3] = dl_detect_out ? proc_dep_vld_vec_24_reg[3] : (proc_24_data_FIFO_blk[3] | proc_24_data_PIPO_blk[3] | proc_24_start_FIFO_blk[3] | proc_24_TLF_FIFO_blk[3] | proc_24_input_sync_blk[3] | proc_24_output_sync_blk[3]);
    assign proc_24_data_FIFO_blk[4] = 1'b0;
    assign proc_24_data_PIPO_blk[4] = 1'b0;
    assign proc_24_start_FIFO_blk[4] = 1'b0;
    assign proc_24_TLF_FIFO_blk[4] = 1'b0;
    assign proc_24_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_24_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_24[4] = dl_detect_out ? proc_dep_vld_vec_24_reg[4] : (proc_24_data_FIFO_blk[4] | proc_24_data_PIPO_blk[4] | proc_24_start_FIFO_blk[4] | proc_24_TLF_FIFO_blk[4] | proc_24_input_sync_blk[4] | proc_24_output_sync_blk[4]);
    assign proc_24_data_FIFO_blk[5] = 1'b0;
    assign proc_24_data_PIPO_blk[5] = 1'b0;
    assign proc_24_start_FIFO_blk[5] = 1'b0;
    assign proc_24_TLF_FIFO_blk[5] = 1'b0;
    assign proc_24_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_24_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_24[5] = dl_detect_out ? proc_dep_vld_vec_24_reg[5] : (proc_24_data_FIFO_blk[5] | proc_24_data_PIPO_blk[5] | proc_24_start_FIFO_blk[5] | proc_24_TLF_FIFO_blk[5] | proc_24_input_sync_blk[5] | proc_24_output_sync_blk[5]);
    assign proc_24_data_FIFO_blk[6] = 1'b0;
    assign proc_24_data_PIPO_blk[6] = 1'b0;
    assign proc_24_start_FIFO_blk[6] = 1'b0;
    assign proc_24_TLF_FIFO_blk[6] = 1'b0;
    assign proc_24_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_24_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_24[6] = dl_detect_out ? proc_dep_vld_vec_24_reg[6] : (proc_24_data_FIFO_blk[6] | proc_24_data_PIPO_blk[6] | proc_24_start_FIFO_blk[6] | proc_24_TLF_FIFO_blk[6] | proc_24_input_sync_blk[6] | proc_24_output_sync_blk[6]);
    assign proc_24_data_FIFO_blk[7] = 1'b0;
    assign proc_24_data_PIPO_blk[7] = 1'b0;
    assign proc_24_start_FIFO_blk[7] = 1'b0;
    assign proc_24_TLF_FIFO_blk[7] = 1'b0;
    assign proc_24_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_24_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_24[7] = dl_detect_out ? proc_dep_vld_vec_24_reg[7] : (proc_24_data_FIFO_blk[7] | proc_24_data_PIPO_blk[7] | proc_24_start_FIFO_blk[7] | proc_24_TLF_FIFO_blk[7] | proc_24_input_sync_blk[7] | proc_24_output_sync_blk[7]);
    assign proc_24_data_FIFO_blk[8] = 1'b0;
    assign proc_24_data_PIPO_blk[8] = 1'b0;
    assign proc_24_start_FIFO_blk[8] = 1'b0;
    assign proc_24_TLF_FIFO_blk[8] = 1'b0;
    assign proc_24_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_24_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_24[8] = dl_detect_out ? proc_dep_vld_vec_24_reg[8] : (proc_24_data_FIFO_blk[8] | proc_24_data_PIPO_blk[8] | proc_24_start_FIFO_blk[8] | proc_24_TLF_FIFO_blk[8] | proc_24_input_sync_blk[8] | proc_24_output_sync_blk[8]);
    assign proc_24_data_FIFO_blk[9] = 1'b0;
    assign proc_24_data_PIPO_blk[9] = 1'b0;
    assign proc_24_start_FIFO_blk[9] = 1'b0;
    assign proc_24_TLF_FIFO_blk[9] = 1'b0;
    assign proc_24_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_24_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_24[9] = dl_detect_out ? proc_dep_vld_vec_24_reg[9] : (proc_24_data_FIFO_blk[9] | proc_24_data_PIPO_blk[9] | proc_24_start_FIFO_blk[9] | proc_24_TLF_FIFO_blk[9] | proc_24_input_sync_blk[9] | proc_24_output_sync_blk[9]);
    assign proc_24_data_FIFO_blk[10] = 1'b0;
    assign proc_24_data_PIPO_blk[10] = 1'b0;
    assign proc_24_start_FIFO_blk[10] = 1'b0;
    assign proc_24_TLF_FIFO_blk[10] = 1'b0;
    assign proc_24_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_24_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_24[10] = dl_detect_out ? proc_dep_vld_vec_24_reg[10] : (proc_24_data_FIFO_blk[10] | proc_24_data_PIPO_blk[10] | proc_24_start_FIFO_blk[10] | proc_24_TLF_FIFO_blk[10] | proc_24_input_sync_blk[10] | proc_24_output_sync_blk[10]);
    assign proc_24_data_FIFO_blk[11] = 1'b0;
    assign proc_24_data_PIPO_blk[11] = 1'b0;
    assign proc_24_start_FIFO_blk[11] = 1'b0;
    assign proc_24_TLF_FIFO_blk[11] = 1'b0;
    assign proc_24_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_24_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_24[11] = dl_detect_out ? proc_dep_vld_vec_24_reg[11] : (proc_24_data_FIFO_blk[11] | proc_24_data_PIPO_blk[11] | proc_24_start_FIFO_blk[11] | proc_24_TLF_FIFO_blk[11] | proc_24_input_sync_blk[11] | proc_24_output_sync_blk[11]);
    assign proc_24_data_FIFO_blk[12] = 1'b0;
    assign proc_24_data_PIPO_blk[12] = 1'b0;
    assign proc_24_start_FIFO_blk[12] = 1'b0;
    assign proc_24_TLF_FIFO_blk[12] = 1'b0;
    assign proc_24_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_24_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_24[12] = dl_detect_out ? proc_dep_vld_vec_24_reg[12] : (proc_24_data_FIFO_blk[12] | proc_24_data_PIPO_blk[12] | proc_24_start_FIFO_blk[12] | proc_24_TLF_FIFO_blk[12] | proc_24_input_sync_blk[12] | proc_24_output_sync_blk[12]);
    assign proc_24_data_FIFO_blk[13] = 1'b0;
    assign proc_24_data_PIPO_blk[13] = 1'b0;
    assign proc_24_start_FIFO_blk[13] = 1'b0;
    assign proc_24_TLF_FIFO_blk[13] = 1'b0;
    assign proc_24_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_24_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_24[13] = dl_detect_out ? proc_dep_vld_vec_24_reg[13] : (proc_24_data_FIFO_blk[13] | proc_24_data_PIPO_blk[13] | proc_24_start_FIFO_blk[13] | proc_24_TLF_FIFO_blk[13] | proc_24_input_sync_blk[13] | proc_24_output_sync_blk[13]);
    assign proc_24_data_FIFO_blk[14] = 1'b0;
    assign proc_24_data_PIPO_blk[14] = 1'b0;
    assign proc_24_start_FIFO_blk[14] = 1'b0;
    assign proc_24_TLF_FIFO_blk[14] = 1'b0;
    assign proc_24_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_24_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_24[14] = dl_detect_out ? proc_dep_vld_vec_24_reg[14] : (proc_24_data_FIFO_blk[14] | proc_24_data_PIPO_blk[14] | proc_24_start_FIFO_blk[14] | proc_24_TLF_FIFO_blk[14] | proc_24_input_sync_blk[14] | proc_24_output_sync_blk[14]);
    assign proc_24_data_FIFO_blk[15] = 1'b0;
    assign proc_24_data_PIPO_blk[15] = 1'b0;
    assign proc_24_start_FIFO_blk[15] = 1'b0;
    assign proc_24_TLF_FIFO_blk[15] = 1'b0;
    assign proc_24_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_24_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_24[15] = dl_detect_out ? proc_dep_vld_vec_24_reg[15] : (proc_24_data_FIFO_blk[15] | proc_24_data_PIPO_blk[15] | proc_24_start_FIFO_blk[15] | proc_24_TLF_FIFO_blk[15] | proc_24_input_sync_blk[15] | proc_24_output_sync_blk[15]);
    assign proc_24_data_FIFO_blk[16] = 1'b0;
    assign proc_24_data_PIPO_blk[16] = 1'b0;
    assign proc_24_start_FIFO_blk[16] = 1'b0;
    assign proc_24_TLF_FIFO_blk[16] = 1'b0;
    assign proc_24_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_24_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_24[16] = dl_detect_out ? proc_dep_vld_vec_24_reg[16] : (proc_24_data_FIFO_blk[16] | proc_24_data_PIPO_blk[16] | proc_24_start_FIFO_blk[16] | proc_24_TLF_FIFO_blk[16] | proc_24_input_sync_blk[16] | proc_24_output_sync_blk[16]);
    assign proc_24_data_FIFO_blk[17] = 1'b0;
    assign proc_24_data_PIPO_blk[17] = 1'b0;
    assign proc_24_start_FIFO_blk[17] = 1'b0;
    assign proc_24_TLF_FIFO_blk[17] = 1'b0;
    assign proc_24_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_24_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_24[17] = dl_detect_out ? proc_dep_vld_vec_24_reg[17] : (proc_24_data_FIFO_blk[17] | proc_24_data_PIPO_blk[17] | proc_24_start_FIFO_blk[17] | proc_24_TLF_FIFO_blk[17] | proc_24_input_sync_blk[17] | proc_24_output_sync_blk[17]);
    assign proc_24_data_FIFO_blk[18] = 1'b0;
    assign proc_24_data_PIPO_blk[18] = 1'b0;
    assign proc_24_start_FIFO_blk[18] = 1'b0;
    assign proc_24_TLF_FIFO_blk[18] = 1'b0;
    assign proc_24_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_24_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_24[18] = dl_detect_out ? proc_dep_vld_vec_24_reg[18] : (proc_24_data_FIFO_blk[18] | proc_24_data_PIPO_blk[18] | proc_24_start_FIFO_blk[18] | proc_24_TLF_FIFO_blk[18] | proc_24_input_sync_blk[18] | proc_24_output_sync_blk[18]);
    assign proc_24_data_FIFO_blk[19] = 1'b0;
    assign proc_24_data_PIPO_blk[19] = 1'b0;
    assign proc_24_start_FIFO_blk[19] = 1'b0;
    assign proc_24_TLF_FIFO_blk[19] = 1'b0;
    assign proc_24_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_24_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_24[19] = dl_detect_out ? proc_dep_vld_vec_24_reg[19] : (proc_24_data_FIFO_blk[19] | proc_24_data_PIPO_blk[19] | proc_24_start_FIFO_blk[19] | proc_24_TLF_FIFO_blk[19] | proc_24_input_sync_blk[19] | proc_24_output_sync_blk[19]);
    assign proc_24_data_FIFO_blk[20] = 1'b0;
    assign proc_24_data_PIPO_blk[20] = 1'b0;
    assign proc_24_start_FIFO_blk[20] = 1'b0;
    assign proc_24_TLF_FIFO_blk[20] = 1'b0;
    assign proc_24_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_24_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_24[20] = dl_detect_out ? proc_dep_vld_vec_24_reg[20] : (proc_24_data_FIFO_blk[20] | proc_24_data_PIPO_blk[20] | proc_24_start_FIFO_blk[20] | proc_24_TLF_FIFO_blk[20] | proc_24_input_sync_blk[20] | proc_24_output_sync_blk[20]);
    assign proc_24_data_FIFO_blk[21] = 1'b0;
    assign proc_24_data_PIPO_blk[21] = 1'b0;
    assign proc_24_start_FIFO_blk[21] = 1'b0;
    assign proc_24_TLF_FIFO_blk[21] = 1'b0;
    assign proc_24_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_24_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_24[21] = dl_detect_out ? proc_dep_vld_vec_24_reg[21] : (proc_24_data_FIFO_blk[21] | proc_24_data_PIPO_blk[21] | proc_24_start_FIFO_blk[21] | proc_24_TLF_FIFO_blk[21] | proc_24_input_sync_blk[21] | proc_24_output_sync_blk[21]);
    assign proc_24_data_FIFO_blk[22] = 1'b0;
    assign proc_24_data_PIPO_blk[22] = 1'b0;
    assign proc_24_start_FIFO_blk[22] = 1'b0;
    assign proc_24_TLF_FIFO_blk[22] = 1'b0;
    assign proc_24_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_24_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_24[22] = dl_detect_out ? proc_dep_vld_vec_24_reg[22] : (proc_24_data_FIFO_blk[22] | proc_24_data_PIPO_blk[22] | proc_24_start_FIFO_blk[22] | proc_24_TLF_FIFO_blk[22] | proc_24_input_sync_blk[22] | proc_24_output_sync_blk[22]);
    assign proc_24_data_FIFO_blk[23] = 1'b0;
    assign proc_24_data_PIPO_blk[23] = 1'b0;
    assign proc_24_start_FIFO_blk[23] = 1'b0;
    assign proc_24_TLF_FIFO_blk[23] = 1'b0;
    assign proc_24_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_24_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_24[23] = dl_detect_out ? proc_dep_vld_vec_24_reg[23] : (proc_24_data_FIFO_blk[23] | proc_24_data_PIPO_blk[23] | proc_24_start_FIFO_blk[23] | proc_24_TLF_FIFO_blk[23] | proc_24_input_sync_blk[23] | proc_24_output_sync_blk[23]);
    assign proc_24_data_FIFO_blk[24] = 1'b0;
    assign proc_24_data_PIPO_blk[24] = 1'b0;
    assign proc_24_start_FIFO_blk[24] = 1'b0;
    assign proc_24_TLF_FIFO_blk[24] = 1'b0;
    assign proc_24_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_24_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_24[24] = dl_detect_out ? proc_dep_vld_vec_24_reg[24] : (proc_24_data_FIFO_blk[24] | proc_24_data_PIPO_blk[24] | proc_24_start_FIFO_blk[24] | proc_24_TLF_FIFO_blk[24] | proc_24_input_sync_blk[24] | proc_24_output_sync_blk[24]);
    assign proc_24_data_FIFO_blk[25] = 1'b0;
    assign proc_24_data_PIPO_blk[25] = 1'b0;
    assign proc_24_start_FIFO_blk[25] = 1'b0;
    assign proc_24_TLF_FIFO_blk[25] = 1'b0;
    assign proc_24_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_24_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_24[25] = dl_detect_out ? proc_dep_vld_vec_24_reg[25] : (proc_24_data_FIFO_blk[25] | proc_24_data_PIPO_blk[25] | proc_24_start_FIFO_blk[25] | proc_24_TLF_FIFO_blk[25] | proc_24_input_sync_blk[25] | proc_24_output_sync_blk[25]);
    assign proc_24_data_FIFO_blk[26] = 1'b0;
    assign proc_24_data_PIPO_blk[26] = 1'b0;
    assign proc_24_start_FIFO_blk[26] = 1'b0;
    assign proc_24_TLF_FIFO_blk[26] = 1'b0;
    assign proc_24_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_24_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_24[26] = dl_detect_out ? proc_dep_vld_vec_24_reg[26] : (proc_24_data_FIFO_blk[26] | proc_24_data_PIPO_blk[26] | proc_24_start_FIFO_blk[26] | proc_24_TLF_FIFO_blk[26] | proc_24_input_sync_blk[26] | proc_24_output_sync_blk[26]);
    assign proc_24_data_FIFO_blk[27] = 1'b0;
    assign proc_24_data_PIPO_blk[27] = 1'b0;
    assign proc_24_start_FIFO_blk[27] = 1'b0;
    assign proc_24_TLF_FIFO_blk[27] = 1'b0;
    assign proc_24_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_24_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_24[27] = dl_detect_out ? proc_dep_vld_vec_24_reg[27] : (proc_24_data_FIFO_blk[27] | proc_24_data_PIPO_blk[27] | proc_24_start_FIFO_blk[27] | proc_24_TLF_FIFO_blk[27] | proc_24_input_sync_blk[27] | proc_24_output_sync_blk[27]);
    assign proc_24_data_FIFO_blk[28] = 1'b0;
    assign proc_24_data_PIPO_blk[28] = 1'b0;
    assign proc_24_start_FIFO_blk[28] = 1'b0;
    assign proc_24_TLF_FIFO_blk[28] = 1'b0;
    assign proc_24_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_24_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_24[28] = dl_detect_out ? proc_dep_vld_vec_24_reg[28] : (proc_24_data_FIFO_blk[28] | proc_24_data_PIPO_blk[28] | proc_24_start_FIFO_blk[28] | proc_24_TLF_FIFO_blk[28] | proc_24_input_sync_blk[28] | proc_24_output_sync_blk[28]);
    assign proc_24_data_FIFO_blk[29] = 1'b0;
    assign proc_24_data_PIPO_blk[29] = 1'b0;
    assign proc_24_start_FIFO_blk[29] = 1'b0;
    assign proc_24_TLF_FIFO_blk[29] = 1'b0;
    assign proc_24_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_24_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_24[29] = dl_detect_out ? proc_dep_vld_vec_24_reg[29] : (proc_24_data_FIFO_blk[29] | proc_24_data_PIPO_blk[29] | proc_24_start_FIFO_blk[29] | proc_24_TLF_FIFO_blk[29] | proc_24_input_sync_blk[29] | proc_24_output_sync_blk[29]);
    assign proc_24_data_FIFO_blk[30] = 1'b0;
    assign proc_24_data_PIPO_blk[30] = 1'b0;
    assign proc_24_start_FIFO_blk[30] = 1'b0;
    assign proc_24_TLF_FIFO_blk[30] = 1'b0;
    assign proc_24_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_24_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_24[30] = dl_detect_out ? proc_dep_vld_vec_24_reg[30] : (proc_24_data_FIFO_blk[30] | proc_24_data_PIPO_blk[30] | proc_24_start_FIFO_blk[30] | proc_24_TLF_FIFO_blk[30] | proc_24_input_sync_blk[30] | proc_24_output_sync_blk[30]);
    assign proc_24_data_FIFO_blk[31] = 1'b0;
    assign proc_24_data_PIPO_blk[31] = 1'b0;
    assign proc_24_start_FIFO_blk[31] = 1'b0;
    assign proc_24_TLF_FIFO_blk[31] = 1'b0;
    assign proc_24_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_24_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_24[31] = dl_detect_out ? proc_dep_vld_vec_24_reg[31] : (proc_24_data_FIFO_blk[31] | proc_24_data_PIPO_blk[31] | proc_24_start_FIFO_blk[31] | proc_24_TLF_FIFO_blk[31] | proc_24_input_sync_blk[31] | proc_24_output_sync_blk[31]);
    assign proc_24_data_FIFO_blk[32] = 1'b0;
    assign proc_24_data_PIPO_blk[32] = 1'b0;
    assign proc_24_start_FIFO_blk[32] = 1'b0;
    assign proc_24_TLF_FIFO_blk[32] = 1'b0;
    assign proc_24_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_19_U0_ap_ready & ProcessingElement_19_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_24_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_24[32] = dl_detect_out ? proc_dep_vld_vec_24_reg[32] : (proc_24_data_FIFO_blk[32] | proc_24_data_PIPO_blk[32] | proc_24_start_FIFO_blk[32] | proc_24_TLF_FIFO_blk[32] | proc_24_input_sync_blk[32] | proc_24_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_24_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_24_reg <= proc_dep_vld_vec_24;
        end
    end
    assign in_chan_dep_vld_vec_24[0] = dep_chan_vld_0_24;
    assign in_chan_dep_data_vec_24[39 : 0] = dep_chan_data_0_24;
    assign token_in_vec_24[0] = token_0_24;
    assign in_chan_dep_vld_vec_24[1] = dep_chan_vld_1_24;
    assign in_chan_dep_data_vec_24[79 : 40] = dep_chan_data_1_24;
    assign token_in_vec_24[1] = token_1_24;
    assign in_chan_dep_vld_vec_24[2] = dep_chan_vld_3_24;
    assign in_chan_dep_data_vec_24[119 : 80] = dep_chan_data_3_24;
    assign token_in_vec_24[2] = token_3_24;
    assign in_chan_dep_vld_vec_24[3] = dep_chan_vld_6_24;
    assign in_chan_dep_data_vec_24[159 : 120] = dep_chan_data_6_24;
    assign token_in_vec_24[3] = token_6_24;
    assign in_chan_dep_vld_vec_24[4] = dep_chan_vld_7_24;
    assign in_chan_dep_data_vec_24[199 : 160] = dep_chan_data_7_24;
    assign token_in_vec_24[4] = token_7_24;
    assign in_chan_dep_vld_vec_24[5] = dep_chan_vld_8_24;
    assign in_chan_dep_data_vec_24[239 : 200] = dep_chan_data_8_24;
    assign token_in_vec_24[5] = token_8_24;
    assign in_chan_dep_vld_vec_24[6] = dep_chan_vld_9_24;
    assign in_chan_dep_data_vec_24[279 : 240] = dep_chan_data_9_24;
    assign token_in_vec_24[6] = token_9_24;
    assign in_chan_dep_vld_vec_24[7] = dep_chan_vld_10_24;
    assign in_chan_dep_data_vec_24[319 : 280] = dep_chan_data_10_24;
    assign token_in_vec_24[7] = token_10_24;
    assign in_chan_dep_vld_vec_24[8] = dep_chan_vld_11_24;
    assign in_chan_dep_data_vec_24[359 : 320] = dep_chan_data_11_24;
    assign token_in_vec_24[8] = token_11_24;
    assign in_chan_dep_vld_vec_24[9] = dep_chan_vld_12_24;
    assign in_chan_dep_data_vec_24[399 : 360] = dep_chan_data_12_24;
    assign token_in_vec_24[9] = token_12_24;
    assign in_chan_dep_vld_vec_24[10] = dep_chan_vld_13_24;
    assign in_chan_dep_data_vec_24[439 : 400] = dep_chan_data_13_24;
    assign token_in_vec_24[10] = token_13_24;
    assign in_chan_dep_vld_vec_24[11] = dep_chan_vld_14_24;
    assign in_chan_dep_data_vec_24[479 : 440] = dep_chan_data_14_24;
    assign token_in_vec_24[11] = token_14_24;
    assign in_chan_dep_vld_vec_24[12] = dep_chan_vld_15_24;
    assign in_chan_dep_data_vec_24[519 : 480] = dep_chan_data_15_24;
    assign token_in_vec_24[12] = token_15_24;
    assign in_chan_dep_vld_vec_24[13] = dep_chan_vld_16_24;
    assign in_chan_dep_data_vec_24[559 : 520] = dep_chan_data_16_24;
    assign token_in_vec_24[13] = token_16_24;
    assign in_chan_dep_vld_vec_24[14] = dep_chan_vld_17_24;
    assign in_chan_dep_data_vec_24[599 : 560] = dep_chan_data_17_24;
    assign token_in_vec_24[14] = token_17_24;
    assign in_chan_dep_vld_vec_24[15] = dep_chan_vld_18_24;
    assign in_chan_dep_data_vec_24[639 : 600] = dep_chan_data_18_24;
    assign token_in_vec_24[15] = token_18_24;
    assign in_chan_dep_vld_vec_24[16] = dep_chan_vld_19_24;
    assign in_chan_dep_data_vec_24[679 : 640] = dep_chan_data_19_24;
    assign token_in_vec_24[16] = token_19_24;
    assign in_chan_dep_vld_vec_24[17] = dep_chan_vld_20_24;
    assign in_chan_dep_data_vec_24[719 : 680] = dep_chan_data_20_24;
    assign token_in_vec_24[17] = token_20_24;
    assign in_chan_dep_vld_vec_24[18] = dep_chan_vld_21_24;
    assign in_chan_dep_data_vec_24[759 : 720] = dep_chan_data_21_24;
    assign token_in_vec_24[18] = token_21_24;
    assign in_chan_dep_vld_vec_24[19] = dep_chan_vld_22_24;
    assign in_chan_dep_data_vec_24[799 : 760] = dep_chan_data_22_24;
    assign token_in_vec_24[19] = token_22_24;
    assign in_chan_dep_vld_vec_24[20] = dep_chan_vld_23_24;
    assign in_chan_dep_data_vec_24[839 : 800] = dep_chan_data_23_24;
    assign token_in_vec_24[20] = token_23_24;
    assign in_chan_dep_vld_vec_24[21] = dep_chan_vld_25_24;
    assign in_chan_dep_data_vec_24[879 : 840] = dep_chan_data_25_24;
    assign token_in_vec_24[21] = token_25_24;
    assign in_chan_dep_vld_vec_24[22] = dep_chan_vld_26_24;
    assign in_chan_dep_data_vec_24[919 : 880] = dep_chan_data_26_24;
    assign token_in_vec_24[22] = token_26_24;
    assign in_chan_dep_vld_vec_24[23] = dep_chan_vld_27_24;
    assign in_chan_dep_data_vec_24[959 : 920] = dep_chan_data_27_24;
    assign token_in_vec_24[23] = token_27_24;
    assign in_chan_dep_vld_vec_24[24] = dep_chan_vld_28_24;
    assign in_chan_dep_data_vec_24[999 : 960] = dep_chan_data_28_24;
    assign token_in_vec_24[24] = token_28_24;
    assign in_chan_dep_vld_vec_24[25] = dep_chan_vld_29_24;
    assign in_chan_dep_data_vec_24[1039 : 1000] = dep_chan_data_29_24;
    assign token_in_vec_24[25] = token_29_24;
    assign in_chan_dep_vld_vec_24[26] = dep_chan_vld_30_24;
    assign in_chan_dep_data_vec_24[1079 : 1040] = dep_chan_data_30_24;
    assign token_in_vec_24[26] = token_30_24;
    assign in_chan_dep_vld_vec_24[27] = dep_chan_vld_31_24;
    assign in_chan_dep_data_vec_24[1119 : 1080] = dep_chan_data_31_24;
    assign token_in_vec_24[27] = token_31_24;
    assign in_chan_dep_vld_vec_24[28] = dep_chan_vld_32_24;
    assign in_chan_dep_data_vec_24[1159 : 1120] = dep_chan_data_32_24;
    assign token_in_vec_24[28] = token_32_24;
    assign in_chan_dep_vld_vec_24[29] = dep_chan_vld_33_24;
    assign in_chan_dep_data_vec_24[1199 : 1160] = dep_chan_data_33_24;
    assign token_in_vec_24[29] = token_33_24;
    assign in_chan_dep_vld_vec_24[30] = dep_chan_vld_34_24;
    assign in_chan_dep_data_vec_24[1239 : 1200] = dep_chan_data_34_24;
    assign token_in_vec_24[30] = token_34_24;
    assign in_chan_dep_vld_vec_24[31] = dep_chan_vld_35_24;
    assign in_chan_dep_data_vec_24[1279 : 1240] = dep_chan_data_35_24;
    assign token_in_vec_24[31] = token_35_24;
    assign in_chan_dep_vld_vec_24[32] = dep_chan_vld_36_24;
    assign in_chan_dep_data_vec_24[1319 : 1280] = dep_chan_data_36_24;
    assign token_in_vec_24[32] = token_36_24;
    assign dep_chan_vld_24_23 = out_chan_dep_vld_vec_24[0];
    assign dep_chan_data_24_23 = out_chan_dep_data_24;
    assign token_24_23 = token_out_vec_24[0];
    assign dep_chan_vld_24_25 = out_chan_dep_vld_vec_24[1];
    assign dep_chan_data_24_25 = out_chan_dep_data_24;
    assign token_24_25 = token_out_vec_24[1];
    assign dep_chan_vld_24_0 = out_chan_dep_vld_vec_24[2];
    assign dep_chan_data_24_0 = out_chan_dep_data_24;
    assign token_24_0 = token_out_vec_24[2];
    assign dep_chan_vld_24_1 = out_chan_dep_vld_vec_24[3];
    assign dep_chan_data_24_1 = out_chan_dep_data_24;
    assign token_24_1 = token_out_vec_24[3];
    assign dep_chan_vld_24_3 = out_chan_dep_vld_vec_24[4];
    assign dep_chan_data_24_3 = out_chan_dep_data_24;
    assign token_24_3 = token_out_vec_24[4];
    assign dep_chan_vld_24_6 = out_chan_dep_vld_vec_24[5];
    assign dep_chan_data_24_6 = out_chan_dep_data_24;
    assign token_24_6 = token_out_vec_24[5];
    assign dep_chan_vld_24_7 = out_chan_dep_vld_vec_24[6];
    assign dep_chan_data_24_7 = out_chan_dep_data_24;
    assign token_24_7 = token_out_vec_24[6];
    assign dep_chan_vld_24_8 = out_chan_dep_vld_vec_24[7];
    assign dep_chan_data_24_8 = out_chan_dep_data_24;
    assign token_24_8 = token_out_vec_24[7];
    assign dep_chan_vld_24_9 = out_chan_dep_vld_vec_24[8];
    assign dep_chan_data_24_9 = out_chan_dep_data_24;
    assign token_24_9 = token_out_vec_24[8];
    assign dep_chan_vld_24_10 = out_chan_dep_vld_vec_24[9];
    assign dep_chan_data_24_10 = out_chan_dep_data_24;
    assign token_24_10 = token_out_vec_24[9];
    assign dep_chan_vld_24_11 = out_chan_dep_vld_vec_24[10];
    assign dep_chan_data_24_11 = out_chan_dep_data_24;
    assign token_24_11 = token_out_vec_24[10];
    assign dep_chan_vld_24_12 = out_chan_dep_vld_vec_24[11];
    assign dep_chan_data_24_12 = out_chan_dep_data_24;
    assign token_24_12 = token_out_vec_24[11];
    assign dep_chan_vld_24_13 = out_chan_dep_vld_vec_24[12];
    assign dep_chan_data_24_13 = out_chan_dep_data_24;
    assign token_24_13 = token_out_vec_24[12];
    assign dep_chan_vld_24_14 = out_chan_dep_vld_vec_24[13];
    assign dep_chan_data_24_14 = out_chan_dep_data_24;
    assign token_24_14 = token_out_vec_24[13];
    assign dep_chan_vld_24_15 = out_chan_dep_vld_vec_24[14];
    assign dep_chan_data_24_15 = out_chan_dep_data_24;
    assign token_24_15 = token_out_vec_24[14];
    assign dep_chan_vld_24_16 = out_chan_dep_vld_vec_24[15];
    assign dep_chan_data_24_16 = out_chan_dep_data_24;
    assign token_24_16 = token_out_vec_24[15];
    assign dep_chan_vld_24_17 = out_chan_dep_vld_vec_24[16];
    assign dep_chan_data_24_17 = out_chan_dep_data_24;
    assign token_24_17 = token_out_vec_24[16];
    assign dep_chan_vld_24_18 = out_chan_dep_vld_vec_24[17];
    assign dep_chan_data_24_18 = out_chan_dep_data_24;
    assign token_24_18 = token_out_vec_24[17];
    assign dep_chan_vld_24_19 = out_chan_dep_vld_vec_24[18];
    assign dep_chan_data_24_19 = out_chan_dep_data_24;
    assign token_24_19 = token_out_vec_24[18];
    assign dep_chan_vld_24_20 = out_chan_dep_vld_vec_24[19];
    assign dep_chan_data_24_20 = out_chan_dep_data_24;
    assign token_24_20 = token_out_vec_24[19];
    assign dep_chan_vld_24_21 = out_chan_dep_vld_vec_24[20];
    assign dep_chan_data_24_21 = out_chan_dep_data_24;
    assign token_24_21 = token_out_vec_24[20];
    assign dep_chan_vld_24_22 = out_chan_dep_vld_vec_24[21];
    assign dep_chan_data_24_22 = out_chan_dep_data_24;
    assign token_24_22 = token_out_vec_24[21];
    assign dep_chan_vld_24_26 = out_chan_dep_vld_vec_24[22];
    assign dep_chan_data_24_26 = out_chan_dep_data_24;
    assign token_24_26 = token_out_vec_24[22];
    assign dep_chan_vld_24_27 = out_chan_dep_vld_vec_24[23];
    assign dep_chan_data_24_27 = out_chan_dep_data_24;
    assign token_24_27 = token_out_vec_24[23];
    assign dep_chan_vld_24_28 = out_chan_dep_vld_vec_24[24];
    assign dep_chan_data_24_28 = out_chan_dep_data_24;
    assign token_24_28 = token_out_vec_24[24];
    assign dep_chan_vld_24_29 = out_chan_dep_vld_vec_24[25];
    assign dep_chan_data_24_29 = out_chan_dep_data_24;
    assign token_24_29 = token_out_vec_24[25];
    assign dep_chan_vld_24_30 = out_chan_dep_vld_vec_24[26];
    assign dep_chan_data_24_30 = out_chan_dep_data_24;
    assign token_24_30 = token_out_vec_24[26];
    assign dep_chan_vld_24_31 = out_chan_dep_vld_vec_24[27];
    assign dep_chan_data_24_31 = out_chan_dep_data_24;
    assign token_24_31 = token_out_vec_24[27];
    assign dep_chan_vld_24_32 = out_chan_dep_vld_vec_24[28];
    assign dep_chan_data_24_32 = out_chan_dep_data_24;
    assign token_24_32 = token_out_vec_24[28];
    assign dep_chan_vld_24_33 = out_chan_dep_vld_vec_24[29];
    assign dep_chan_data_24_33 = out_chan_dep_data_24;
    assign token_24_33 = token_out_vec_24[29];
    assign dep_chan_vld_24_34 = out_chan_dep_vld_vec_24[30];
    assign dep_chan_data_24_34 = out_chan_dep_data_24;
    assign token_24_34 = token_out_vec_24[30];
    assign dep_chan_vld_24_35 = out_chan_dep_vld_vec_24[31];
    assign dep_chan_data_24_35 = out_chan_dep_data_24;
    assign token_24_35 = token_out_vec_24[31];
    assign dep_chan_vld_24_36 = out_chan_dep_vld_vec_24[32];
    assign dep_chan_data_24_36 = out_chan_dep_data_24;
    assign token_24_36 = token_out_vec_24[32];

    // Process: ProcessingElement_20_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 25, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_25 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_25),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_25),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_25),
        .token_in_vec(token_in_vec_25),
        .dl_detect_in(dl_detect_out),
        .origin(origin[25]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_25),
        .out_chan_dep_data(out_chan_dep_data_25),
        .token_out_vec(token_out_vec_25),
        .dl_detect_out(dl_in_vec[25]));

    assign proc_25_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_19_blk_n) | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_19_blk_n) | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_WriteC_Flattened_fu_179.cPipes_19_blk_n);
    assign proc_25_data_PIPO_blk[0] = 1'b0;
    assign proc_25_start_FIFO_blk[0] = 1'b0;
    assign proc_25_TLF_FIFO_blk[0] = 1'b0;
    assign proc_25_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_25_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_25[0] = dl_detect_out ? proc_dep_vld_vec_25_reg[0] : (proc_25_data_FIFO_blk[0] | proc_25_data_PIPO_blk[0] | proc_25_start_FIFO_blk[0] | proc_25_TLF_FIFO_blk[0] | proc_25_input_sync_blk[0] | proc_25_output_sync_blk[0]);
    assign proc_25_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_20_blk_n) | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_20_blk_n) | (~ProcessingElement_20_U0.grp_ProcessingElement_20_Pipeline_WriteC_Flattened_fu_179.cPipes_20_blk_n);
    assign proc_25_data_PIPO_blk[1] = 1'b0;
    assign proc_25_start_FIFO_blk[1] = 1'b0;
    assign proc_25_TLF_FIFO_blk[1] = 1'b0;
    assign proc_25_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_25_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_25[1] = dl_detect_out ? proc_dep_vld_vec_25_reg[1] : (proc_25_data_FIFO_blk[1] | proc_25_data_PIPO_blk[1] | proc_25_start_FIFO_blk[1] | proc_25_TLF_FIFO_blk[1] | proc_25_input_sync_blk[1] | proc_25_output_sync_blk[1]);
    assign proc_25_data_FIFO_blk[2] = 1'b0;
    assign proc_25_data_PIPO_blk[2] = 1'b0;
    assign proc_25_start_FIFO_blk[2] = 1'b0;
    assign proc_25_TLF_FIFO_blk[2] = 1'b0;
    assign proc_25_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_25_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_25[2] = dl_detect_out ? proc_dep_vld_vec_25_reg[2] : (proc_25_data_FIFO_blk[2] | proc_25_data_PIPO_blk[2] | proc_25_start_FIFO_blk[2] | proc_25_TLF_FIFO_blk[2] | proc_25_input_sync_blk[2] | proc_25_output_sync_blk[2]);
    assign proc_25_data_FIFO_blk[3] = 1'b0;
    assign proc_25_data_PIPO_blk[3] = 1'b0;
    assign proc_25_start_FIFO_blk[3] = 1'b0;
    assign proc_25_TLF_FIFO_blk[3] = 1'b0;
    assign proc_25_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_25_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_25[3] = dl_detect_out ? proc_dep_vld_vec_25_reg[3] : (proc_25_data_FIFO_blk[3] | proc_25_data_PIPO_blk[3] | proc_25_start_FIFO_blk[3] | proc_25_TLF_FIFO_blk[3] | proc_25_input_sync_blk[3] | proc_25_output_sync_blk[3]);
    assign proc_25_data_FIFO_blk[4] = 1'b0;
    assign proc_25_data_PIPO_blk[4] = 1'b0;
    assign proc_25_start_FIFO_blk[4] = 1'b0;
    assign proc_25_TLF_FIFO_blk[4] = 1'b0;
    assign proc_25_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_25_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_25[4] = dl_detect_out ? proc_dep_vld_vec_25_reg[4] : (proc_25_data_FIFO_blk[4] | proc_25_data_PIPO_blk[4] | proc_25_start_FIFO_blk[4] | proc_25_TLF_FIFO_blk[4] | proc_25_input_sync_blk[4] | proc_25_output_sync_blk[4]);
    assign proc_25_data_FIFO_blk[5] = 1'b0;
    assign proc_25_data_PIPO_blk[5] = 1'b0;
    assign proc_25_start_FIFO_blk[5] = 1'b0;
    assign proc_25_TLF_FIFO_blk[5] = 1'b0;
    assign proc_25_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_25_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_25[5] = dl_detect_out ? proc_dep_vld_vec_25_reg[5] : (proc_25_data_FIFO_blk[5] | proc_25_data_PIPO_blk[5] | proc_25_start_FIFO_blk[5] | proc_25_TLF_FIFO_blk[5] | proc_25_input_sync_blk[5] | proc_25_output_sync_blk[5]);
    assign proc_25_data_FIFO_blk[6] = 1'b0;
    assign proc_25_data_PIPO_blk[6] = 1'b0;
    assign proc_25_start_FIFO_blk[6] = 1'b0;
    assign proc_25_TLF_FIFO_blk[6] = 1'b0;
    assign proc_25_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_25_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_25[6] = dl_detect_out ? proc_dep_vld_vec_25_reg[6] : (proc_25_data_FIFO_blk[6] | proc_25_data_PIPO_blk[6] | proc_25_start_FIFO_blk[6] | proc_25_TLF_FIFO_blk[6] | proc_25_input_sync_blk[6] | proc_25_output_sync_blk[6]);
    assign proc_25_data_FIFO_blk[7] = 1'b0;
    assign proc_25_data_PIPO_blk[7] = 1'b0;
    assign proc_25_start_FIFO_blk[7] = 1'b0;
    assign proc_25_TLF_FIFO_blk[7] = 1'b0;
    assign proc_25_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_25_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_25[7] = dl_detect_out ? proc_dep_vld_vec_25_reg[7] : (proc_25_data_FIFO_blk[7] | proc_25_data_PIPO_blk[7] | proc_25_start_FIFO_blk[7] | proc_25_TLF_FIFO_blk[7] | proc_25_input_sync_blk[7] | proc_25_output_sync_blk[7]);
    assign proc_25_data_FIFO_blk[8] = 1'b0;
    assign proc_25_data_PIPO_blk[8] = 1'b0;
    assign proc_25_start_FIFO_blk[8] = 1'b0;
    assign proc_25_TLF_FIFO_blk[8] = 1'b0;
    assign proc_25_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_25_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_25[8] = dl_detect_out ? proc_dep_vld_vec_25_reg[8] : (proc_25_data_FIFO_blk[8] | proc_25_data_PIPO_blk[8] | proc_25_start_FIFO_blk[8] | proc_25_TLF_FIFO_blk[8] | proc_25_input_sync_blk[8] | proc_25_output_sync_blk[8]);
    assign proc_25_data_FIFO_blk[9] = 1'b0;
    assign proc_25_data_PIPO_blk[9] = 1'b0;
    assign proc_25_start_FIFO_blk[9] = 1'b0;
    assign proc_25_TLF_FIFO_blk[9] = 1'b0;
    assign proc_25_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_25_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_25[9] = dl_detect_out ? proc_dep_vld_vec_25_reg[9] : (proc_25_data_FIFO_blk[9] | proc_25_data_PIPO_blk[9] | proc_25_start_FIFO_blk[9] | proc_25_TLF_FIFO_blk[9] | proc_25_input_sync_blk[9] | proc_25_output_sync_blk[9]);
    assign proc_25_data_FIFO_blk[10] = 1'b0;
    assign proc_25_data_PIPO_blk[10] = 1'b0;
    assign proc_25_start_FIFO_blk[10] = 1'b0;
    assign proc_25_TLF_FIFO_blk[10] = 1'b0;
    assign proc_25_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_25_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_25[10] = dl_detect_out ? proc_dep_vld_vec_25_reg[10] : (proc_25_data_FIFO_blk[10] | proc_25_data_PIPO_blk[10] | proc_25_start_FIFO_blk[10] | proc_25_TLF_FIFO_blk[10] | proc_25_input_sync_blk[10] | proc_25_output_sync_blk[10]);
    assign proc_25_data_FIFO_blk[11] = 1'b0;
    assign proc_25_data_PIPO_blk[11] = 1'b0;
    assign proc_25_start_FIFO_blk[11] = 1'b0;
    assign proc_25_TLF_FIFO_blk[11] = 1'b0;
    assign proc_25_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_25_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_25[11] = dl_detect_out ? proc_dep_vld_vec_25_reg[11] : (proc_25_data_FIFO_blk[11] | proc_25_data_PIPO_blk[11] | proc_25_start_FIFO_blk[11] | proc_25_TLF_FIFO_blk[11] | proc_25_input_sync_blk[11] | proc_25_output_sync_blk[11]);
    assign proc_25_data_FIFO_blk[12] = 1'b0;
    assign proc_25_data_PIPO_blk[12] = 1'b0;
    assign proc_25_start_FIFO_blk[12] = 1'b0;
    assign proc_25_TLF_FIFO_blk[12] = 1'b0;
    assign proc_25_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_25_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_25[12] = dl_detect_out ? proc_dep_vld_vec_25_reg[12] : (proc_25_data_FIFO_blk[12] | proc_25_data_PIPO_blk[12] | proc_25_start_FIFO_blk[12] | proc_25_TLF_FIFO_blk[12] | proc_25_input_sync_blk[12] | proc_25_output_sync_blk[12]);
    assign proc_25_data_FIFO_blk[13] = 1'b0;
    assign proc_25_data_PIPO_blk[13] = 1'b0;
    assign proc_25_start_FIFO_blk[13] = 1'b0;
    assign proc_25_TLF_FIFO_blk[13] = 1'b0;
    assign proc_25_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_25_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_25[13] = dl_detect_out ? proc_dep_vld_vec_25_reg[13] : (proc_25_data_FIFO_blk[13] | proc_25_data_PIPO_blk[13] | proc_25_start_FIFO_blk[13] | proc_25_TLF_FIFO_blk[13] | proc_25_input_sync_blk[13] | proc_25_output_sync_blk[13]);
    assign proc_25_data_FIFO_blk[14] = 1'b0;
    assign proc_25_data_PIPO_blk[14] = 1'b0;
    assign proc_25_start_FIFO_blk[14] = 1'b0;
    assign proc_25_TLF_FIFO_blk[14] = 1'b0;
    assign proc_25_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_25_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_25[14] = dl_detect_out ? proc_dep_vld_vec_25_reg[14] : (proc_25_data_FIFO_blk[14] | proc_25_data_PIPO_blk[14] | proc_25_start_FIFO_blk[14] | proc_25_TLF_FIFO_blk[14] | proc_25_input_sync_blk[14] | proc_25_output_sync_blk[14]);
    assign proc_25_data_FIFO_blk[15] = 1'b0;
    assign proc_25_data_PIPO_blk[15] = 1'b0;
    assign proc_25_start_FIFO_blk[15] = 1'b0;
    assign proc_25_TLF_FIFO_blk[15] = 1'b0;
    assign proc_25_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_25_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_25[15] = dl_detect_out ? proc_dep_vld_vec_25_reg[15] : (proc_25_data_FIFO_blk[15] | proc_25_data_PIPO_blk[15] | proc_25_start_FIFO_blk[15] | proc_25_TLF_FIFO_blk[15] | proc_25_input_sync_blk[15] | proc_25_output_sync_blk[15]);
    assign proc_25_data_FIFO_blk[16] = 1'b0;
    assign proc_25_data_PIPO_blk[16] = 1'b0;
    assign proc_25_start_FIFO_blk[16] = 1'b0;
    assign proc_25_TLF_FIFO_blk[16] = 1'b0;
    assign proc_25_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_25_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_25[16] = dl_detect_out ? proc_dep_vld_vec_25_reg[16] : (proc_25_data_FIFO_blk[16] | proc_25_data_PIPO_blk[16] | proc_25_start_FIFO_blk[16] | proc_25_TLF_FIFO_blk[16] | proc_25_input_sync_blk[16] | proc_25_output_sync_blk[16]);
    assign proc_25_data_FIFO_blk[17] = 1'b0;
    assign proc_25_data_PIPO_blk[17] = 1'b0;
    assign proc_25_start_FIFO_blk[17] = 1'b0;
    assign proc_25_TLF_FIFO_blk[17] = 1'b0;
    assign proc_25_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_25_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_25[17] = dl_detect_out ? proc_dep_vld_vec_25_reg[17] : (proc_25_data_FIFO_blk[17] | proc_25_data_PIPO_blk[17] | proc_25_start_FIFO_blk[17] | proc_25_TLF_FIFO_blk[17] | proc_25_input_sync_blk[17] | proc_25_output_sync_blk[17]);
    assign proc_25_data_FIFO_blk[18] = 1'b0;
    assign proc_25_data_PIPO_blk[18] = 1'b0;
    assign proc_25_start_FIFO_blk[18] = 1'b0;
    assign proc_25_TLF_FIFO_blk[18] = 1'b0;
    assign proc_25_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_25_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_25[18] = dl_detect_out ? proc_dep_vld_vec_25_reg[18] : (proc_25_data_FIFO_blk[18] | proc_25_data_PIPO_blk[18] | proc_25_start_FIFO_blk[18] | proc_25_TLF_FIFO_blk[18] | proc_25_input_sync_blk[18] | proc_25_output_sync_blk[18]);
    assign proc_25_data_FIFO_blk[19] = 1'b0;
    assign proc_25_data_PIPO_blk[19] = 1'b0;
    assign proc_25_start_FIFO_blk[19] = 1'b0;
    assign proc_25_TLF_FIFO_blk[19] = 1'b0;
    assign proc_25_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_25_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_25[19] = dl_detect_out ? proc_dep_vld_vec_25_reg[19] : (proc_25_data_FIFO_blk[19] | proc_25_data_PIPO_blk[19] | proc_25_start_FIFO_blk[19] | proc_25_TLF_FIFO_blk[19] | proc_25_input_sync_blk[19] | proc_25_output_sync_blk[19]);
    assign proc_25_data_FIFO_blk[20] = 1'b0;
    assign proc_25_data_PIPO_blk[20] = 1'b0;
    assign proc_25_start_FIFO_blk[20] = 1'b0;
    assign proc_25_TLF_FIFO_blk[20] = 1'b0;
    assign proc_25_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_25_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_25[20] = dl_detect_out ? proc_dep_vld_vec_25_reg[20] : (proc_25_data_FIFO_blk[20] | proc_25_data_PIPO_blk[20] | proc_25_start_FIFO_blk[20] | proc_25_TLF_FIFO_blk[20] | proc_25_input_sync_blk[20] | proc_25_output_sync_blk[20]);
    assign proc_25_data_FIFO_blk[21] = 1'b0;
    assign proc_25_data_PIPO_blk[21] = 1'b0;
    assign proc_25_start_FIFO_blk[21] = 1'b0;
    assign proc_25_TLF_FIFO_blk[21] = 1'b0;
    assign proc_25_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_25_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_25[21] = dl_detect_out ? proc_dep_vld_vec_25_reg[21] : (proc_25_data_FIFO_blk[21] | proc_25_data_PIPO_blk[21] | proc_25_start_FIFO_blk[21] | proc_25_TLF_FIFO_blk[21] | proc_25_input_sync_blk[21] | proc_25_output_sync_blk[21]);
    assign proc_25_data_FIFO_blk[22] = 1'b0;
    assign proc_25_data_PIPO_blk[22] = 1'b0;
    assign proc_25_start_FIFO_blk[22] = 1'b0;
    assign proc_25_TLF_FIFO_blk[22] = 1'b0;
    assign proc_25_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_25_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_25[22] = dl_detect_out ? proc_dep_vld_vec_25_reg[22] : (proc_25_data_FIFO_blk[22] | proc_25_data_PIPO_blk[22] | proc_25_start_FIFO_blk[22] | proc_25_TLF_FIFO_blk[22] | proc_25_input_sync_blk[22] | proc_25_output_sync_blk[22]);
    assign proc_25_data_FIFO_blk[23] = 1'b0;
    assign proc_25_data_PIPO_blk[23] = 1'b0;
    assign proc_25_start_FIFO_blk[23] = 1'b0;
    assign proc_25_TLF_FIFO_blk[23] = 1'b0;
    assign proc_25_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_25_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_25[23] = dl_detect_out ? proc_dep_vld_vec_25_reg[23] : (proc_25_data_FIFO_blk[23] | proc_25_data_PIPO_blk[23] | proc_25_start_FIFO_blk[23] | proc_25_TLF_FIFO_blk[23] | proc_25_input_sync_blk[23] | proc_25_output_sync_blk[23]);
    assign proc_25_data_FIFO_blk[24] = 1'b0;
    assign proc_25_data_PIPO_blk[24] = 1'b0;
    assign proc_25_start_FIFO_blk[24] = 1'b0;
    assign proc_25_TLF_FIFO_blk[24] = 1'b0;
    assign proc_25_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_25_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_25[24] = dl_detect_out ? proc_dep_vld_vec_25_reg[24] : (proc_25_data_FIFO_blk[24] | proc_25_data_PIPO_blk[24] | proc_25_start_FIFO_blk[24] | proc_25_TLF_FIFO_blk[24] | proc_25_input_sync_blk[24] | proc_25_output_sync_blk[24]);
    assign proc_25_data_FIFO_blk[25] = 1'b0;
    assign proc_25_data_PIPO_blk[25] = 1'b0;
    assign proc_25_start_FIFO_blk[25] = 1'b0;
    assign proc_25_TLF_FIFO_blk[25] = 1'b0;
    assign proc_25_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_25_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_25[25] = dl_detect_out ? proc_dep_vld_vec_25_reg[25] : (proc_25_data_FIFO_blk[25] | proc_25_data_PIPO_blk[25] | proc_25_start_FIFO_blk[25] | proc_25_TLF_FIFO_blk[25] | proc_25_input_sync_blk[25] | proc_25_output_sync_blk[25]);
    assign proc_25_data_FIFO_blk[26] = 1'b0;
    assign proc_25_data_PIPO_blk[26] = 1'b0;
    assign proc_25_start_FIFO_blk[26] = 1'b0;
    assign proc_25_TLF_FIFO_blk[26] = 1'b0;
    assign proc_25_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_25_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_25[26] = dl_detect_out ? proc_dep_vld_vec_25_reg[26] : (proc_25_data_FIFO_blk[26] | proc_25_data_PIPO_blk[26] | proc_25_start_FIFO_blk[26] | proc_25_TLF_FIFO_blk[26] | proc_25_input_sync_blk[26] | proc_25_output_sync_blk[26]);
    assign proc_25_data_FIFO_blk[27] = 1'b0;
    assign proc_25_data_PIPO_blk[27] = 1'b0;
    assign proc_25_start_FIFO_blk[27] = 1'b0;
    assign proc_25_TLF_FIFO_blk[27] = 1'b0;
    assign proc_25_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_25_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_25[27] = dl_detect_out ? proc_dep_vld_vec_25_reg[27] : (proc_25_data_FIFO_blk[27] | proc_25_data_PIPO_blk[27] | proc_25_start_FIFO_blk[27] | proc_25_TLF_FIFO_blk[27] | proc_25_input_sync_blk[27] | proc_25_output_sync_blk[27]);
    assign proc_25_data_FIFO_blk[28] = 1'b0;
    assign proc_25_data_PIPO_blk[28] = 1'b0;
    assign proc_25_start_FIFO_blk[28] = 1'b0;
    assign proc_25_TLF_FIFO_blk[28] = 1'b0;
    assign proc_25_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_25_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_25[28] = dl_detect_out ? proc_dep_vld_vec_25_reg[28] : (proc_25_data_FIFO_blk[28] | proc_25_data_PIPO_blk[28] | proc_25_start_FIFO_blk[28] | proc_25_TLF_FIFO_blk[28] | proc_25_input_sync_blk[28] | proc_25_output_sync_blk[28]);
    assign proc_25_data_FIFO_blk[29] = 1'b0;
    assign proc_25_data_PIPO_blk[29] = 1'b0;
    assign proc_25_start_FIFO_blk[29] = 1'b0;
    assign proc_25_TLF_FIFO_blk[29] = 1'b0;
    assign proc_25_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_25_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_25[29] = dl_detect_out ? proc_dep_vld_vec_25_reg[29] : (proc_25_data_FIFO_blk[29] | proc_25_data_PIPO_blk[29] | proc_25_start_FIFO_blk[29] | proc_25_TLF_FIFO_blk[29] | proc_25_input_sync_blk[29] | proc_25_output_sync_blk[29]);
    assign proc_25_data_FIFO_blk[30] = 1'b0;
    assign proc_25_data_PIPO_blk[30] = 1'b0;
    assign proc_25_start_FIFO_blk[30] = 1'b0;
    assign proc_25_TLF_FIFO_blk[30] = 1'b0;
    assign proc_25_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_25_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_25[30] = dl_detect_out ? proc_dep_vld_vec_25_reg[30] : (proc_25_data_FIFO_blk[30] | proc_25_data_PIPO_blk[30] | proc_25_start_FIFO_blk[30] | proc_25_TLF_FIFO_blk[30] | proc_25_input_sync_blk[30] | proc_25_output_sync_blk[30]);
    assign proc_25_data_FIFO_blk[31] = 1'b0;
    assign proc_25_data_PIPO_blk[31] = 1'b0;
    assign proc_25_start_FIFO_blk[31] = 1'b0;
    assign proc_25_TLF_FIFO_blk[31] = 1'b0;
    assign proc_25_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_25_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_25[31] = dl_detect_out ? proc_dep_vld_vec_25_reg[31] : (proc_25_data_FIFO_blk[31] | proc_25_data_PIPO_blk[31] | proc_25_start_FIFO_blk[31] | proc_25_TLF_FIFO_blk[31] | proc_25_input_sync_blk[31] | proc_25_output_sync_blk[31]);
    assign proc_25_data_FIFO_blk[32] = 1'b0;
    assign proc_25_data_PIPO_blk[32] = 1'b0;
    assign proc_25_start_FIFO_blk[32] = 1'b0;
    assign proc_25_TLF_FIFO_blk[32] = 1'b0;
    assign proc_25_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_20_U0_ap_ready & ProcessingElement_20_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_25_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_25[32] = dl_detect_out ? proc_dep_vld_vec_25_reg[32] : (proc_25_data_FIFO_blk[32] | proc_25_data_PIPO_blk[32] | proc_25_start_FIFO_blk[32] | proc_25_TLF_FIFO_blk[32] | proc_25_input_sync_blk[32] | proc_25_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_25_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_25_reg <= proc_dep_vld_vec_25;
        end
    end
    assign in_chan_dep_vld_vec_25[0] = dep_chan_vld_0_25;
    assign in_chan_dep_data_vec_25[39 : 0] = dep_chan_data_0_25;
    assign token_in_vec_25[0] = token_0_25;
    assign in_chan_dep_vld_vec_25[1] = dep_chan_vld_1_25;
    assign in_chan_dep_data_vec_25[79 : 40] = dep_chan_data_1_25;
    assign token_in_vec_25[1] = token_1_25;
    assign in_chan_dep_vld_vec_25[2] = dep_chan_vld_3_25;
    assign in_chan_dep_data_vec_25[119 : 80] = dep_chan_data_3_25;
    assign token_in_vec_25[2] = token_3_25;
    assign in_chan_dep_vld_vec_25[3] = dep_chan_vld_6_25;
    assign in_chan_dep_data_vec_25[159 : 120] = dep_chan_data_6_25;
    assign token_in_vec_25[3] = token_6_25;
    assign in_chan_dep_vld_vec_25[4] = dep_chan_vld_7_25;
    assign in_chan_dep_data_vec_25[199 : 160] = dep_chan_data_7_25;
    assign token_in_vec_25[4] = token_7_25;
    assign in_chan_dep_vld_vec_25[5] = dep_chan_vld_8_25;
    assign in_chan_dep_data_vec_25[239 : 200] = dep_chan_data_8_25;
    assign token_in_vec_25[5] = token_8_25;
    assign in_chan_dep_vld_vec_25[6] = dep_chan_vld_9_25;
    assign in_chan_dep_data_vec_25[279 : 240] = dep_chan_data_9_25;
    assign token_in_vec_25[6] = token_9_25;
    assign in_chan_dep_vld_vec_25[7] = dep_chan_vld_10_25;
    assign in_chan_dep_data_vec_25[319 : 280] = dep_chan_data_10_25;
    assign token_in_vec_25[7] = token_10_25;
    assign in_chan_dep_vld_vec_25[8] = dep_chan_vld_11_25;
    assign in_chan_dep_data_vec_25[359 : 320] = dep_chan_data_11_25;
    assign token_in_vec_25[8] = token_11_25;
    assign in_chan_dep_vld_vec_25[9] = dep_chan_vld_12_25;
    assign in_chan_dep_data_vec_25[399 : 360] = dep_chan_data_12_25;
    assign token_in_vec_25[9] = token_12_25;
    assign in_chan_dep_vld_vec_25[10] = dep_chan_vld_13_25;
    assign in_chan_dep_data_vec_25[439 : 400] = dep_chan_data_13_25;
    assign token_in_vec_25[10] = token_13_25;
    assign in_chan_dep_vld_vec_25[11] = dep_chan_vld_14_25;
    assign in_chan_dep_data_vec_25[479 : 440] = dep_chan_data_14_25;
    assign token_in_vec_25[11] = token_14_25;
    assign in_chan_dep_vld_vec_25[12] = dep_chan_vld_15_25;
    assign in_chan_dep_data_vec_25[519 : 480] = dep_chan_data_15_25;
    assign token_in_vec_25[12] = token_15_25;
    assign in_chan_dep_vld_vec_25[13] = dep_chan_vld_16_25;
    assign in_chan_dep_data_vec_25[559 : 520] = dep_chan_data_16_25;
    assign token_in_vec_25[13] = token_16_25;
    assign in_chan_dep_vld_vec_25[14] = dep_chan_vld_17_25;
    assign in_chan_dep_data_vec_25[599 : 560] = dep_chan_data_17_25;
    assign token_in_vec_25[14] = token_17_25;
    assign in_chan_dep_vld_vec_25[15] = dep_chan_vld_18_25;
    assign in_chan_dep_data_vec_25[639 : 600] = dep_chan_data_18_25;
    assign token_in_vec_25[15] = token_18_25;
    assign in_chan_dep_vld_vec_25[16] = dep_chan_vld_19_25;
    assign in_chan_dep_data_vec_25[679 : 640] = dep_chan_data_19_25;
    assign token_in_vec_25[16] = token_19_25;
    assign in_chan_dep_vld_vec_25[17] = dep_chan_vld_20_25;
    assign in_chan_dep_data_vec_25[719 : 680] = dep_chan_data_20_25;
    assign token_in_vec_25[17] = token_20_25;
    assign in_chan_dep_vld_vec_25[18] = dep_chan_vld_21_25;
    assign in_chan_dep_data_vec_25[759 : 720] = dep_chan_data_21_25;
    assign token_in_vec_25[18] = token_21_25;
    assign in_chan_dep_vld_vec_25[19] = dep_chan_vld_22_25;
    assign in_chan_dep_data_vec_25[799 : 760] = dep_chan_data_22_25;
    assign token_in_vec_25[19] = token_22_25;
    assign in_chan_dep_vld_vec_25[20] = dep_chan_vld_23_25;
    assign in_chan_dep_data_vec_25[839 : 800] = dep_chan_data_23_25;
    assign token_in_vec_25[20] = token_23_25;
    assign in_chan_dep_vld_vec_25[21] = dep_chan_vld_24_25;
    assign in_chan_dep_data_vec_25[879 : 840] = dep_chan_data_24_25;
    assign token_in_vec_25[21] = token_24_25;
    assign in_chan_dep_vld_vec_25[22] = dep_chan_vld_26_25;
    assign in_chan_dep_data_vec_25[919 : 880] = dep_chan_data_26_25;
    assign token_in_vec_25[22] = token_26_25;
    assign in_chan_dep_vld_vec_25[23] = dep_chan_vld_27_25;
    assign in_chan_dep_data_vec_25[959 : 920] = dep_chan_data_27_25;
    assign token_in_vec_25[23] = token_27_25;
    assign in_chan_dep_vld_vec_25[24] = dep_chan_vld_28_25;
    assign in_chan_dep_data_vec_25[999 : 960] = dep_chan_data_28_25;
    assign token_in_vec_25[24] = token_28_25;
    assign in_chan_dep_vld_vec_25[25] = dep_chan_vld_29_25;
    assign in_chan_dep_data_vec_25[1039 : 1000] = dep_chan_data_29_25;
    assign token_in_vec_25[25] = token_29_25;
    assign in_chan_dep_vld_vec_25[26] = dep_chan_vld_30_25;
    assign in_chan_dep_data_vec_25[1079 : 1040] = dep_chan_data_30_25;
    assign token_in_vec_25[26] = token_30_25;
    assign in_chan_dep_vld_vec_25[27] = dep_chan_vld_31_25;
    assign in_chan_dep_data_vec_25[1119 : 1080] = dep_chan_data_31_25;
    assign token_in_vec_25[27] = token_31_25;
    assign in_chan_dep_vld_vec_25[28] = dep_chan_vld_32_25;
    assign in_chan_dep_data_vec_25[1159 : 1120] = dep_chan_data_32_25;
    assign token_in_vec_25[28] = token_32_25;
    assign in_chan_dep_vld_vec_25[29] = dep_chan_vld_33_25;
    assign in_chan_dep_data_vec_25[1199 : 1160] = dep_chan_data_33_25;
    assign token_in_vec_25[29] = token_33_25;
    assign in_chan_dep_vld_vec_25[30] = dep_chan_vld_34_25;
    assign in_chan_dep_data_vec_25[1239 : 1200] = dep_chan_data_34_25;
    assign token_in_vec_25[30] = token_34_25;
    assign in_chan_dep_vld_vec_25[31] = dep_chan_vld_35_25;
    assign in_chan_dep_data_vec_25[1279 : 1240] = dep_chan_data_35_25;
    assign token_in_vec_25[31] = token_35_25;
    assign in_chan_dep_vld_vec_25[32] = dep_chan_vld_36_25;
    assign in_chan_dep_data_vec_25[1319 : 1280] = dep_chan_data_36_25;
    assign token_in_vec_25[32] = token_36_25;
    assign dep_chan_vld_25_24 = out_chan_dep_vld_vec_25[0];
    assign dep_chan_data_25_24 = out_chan_dep_data_25;
    assign token_25_24 = token_out_vec_25[0];
    assign dep_chan_vld_25_26 = out_chan_dep_vld_vec_25[1];
    assign dep_chan_data_25_26 = out_chan_dep_data_25;
    assign token_25_26 = token_out_vec_25[1];
    assign dep_chan_vld_25_0 = out_chan_dep_vld_vec_25[2];
    assign dep_chan_data_25_0 = out_chan_dep_data_25;
    assign token_25_0 = token_out_vec_25[2];
    assign dep_chan_vld_25_1 = out_chan_dep_vld_vec_25[3];
    assign dep_chan_data_25_1 = out_chan_dep_data_25;
    assign token_25_1 = token_out_vec_25[3];
    assign dep_chan_vld_25_3 = out_chan_dep_vld_vec_25[4];
    assign dep_chan_data_25_3 = out_chan_dep_data_25;
    assign token_25_3 = token_out_vec_25[4];
    assign dep_chan_vld_25_6 = out_chan_dep_vld_vec_25[5];
    assign dep_chan_data_25_6 = out_chan_dep_data_25;
    assign token_25_6 = token_out_vec_25[5];
    assign dep_chan_vld_25_7 = out_chan_dep_vld_vec_25[6];
    assign dep_chan_data_25_7 = out_chan_dep_data_25;
    assign token_25_7 = token_out_vec_25[6];
    assign dep_chan_vld_25_8 = out_chan_dep_vld_vec_25[7];
    assign dep_chan_data_25_8 = out_chan_dep_data_25;
    assign token_25_8 = token_out_vec_25[7];
    assign dep_chan_vld_25_9 = out_chan_dep_vld_vec_25[8];
    assign dep_chan_data_25_9 = out_chan_dep_data_25;
    assign token_25_9 = token_out_vec_25[8];
    assign dep_chan_vld_25_10 = out_chan_dep_vld_vec_25[9];
    assign dep_chan_data_25_10 = out_chan_dep_data_25;
    assign token_25_10 = token_out_vec_25[9];
    assign dep_chan_vld_25_11 = out_chan_dep_vld_vec_25[10];
    assign dep_chan_data_25_11 = out_chan_dep_data_25;
    assign token_25_11 = token_out_vec_25[10];
    assign dep_chan_vld_25_12 = out_chan_dep_vld_vec_25[11];
    assign dep_chan_data_25_12 = out_chan_dep_data_25;
    assign token_25_12 = token_out_vec_25[11];
    assign dep_chan_vld_25_13 = out_chan_dep_vld_vec_25[12];
    assign dep_chan_data_25_13 = out_chan_dep_data_25;
    assign token_25_13 = token_out_vec_25[12];
    assign dep_chan_vld_25_14 = out_chan_dep_vld_vec_25[13];
    assign dep_chan_data_25_14 = out_chan_dep_data_25;
    assign token_25_14 = token_out_vec_25[13];
    assign dep_chan_vld_25_15 = out_chan_dep_vld_vec_25[14];
    assign dep_chan_data_25_15 = out_chan_dep_data_25;
    assign token_25_15 = token_out_vec_25[14];
    assign dep_chan_vld_25_16 = out_chan_dep_vld_vec_25[15];
    assign dep_chan_data_25_16 = out_chan_dep_data_25;
    assign token_25_16 = token_out_vec_25[15];
    assign dep_chan_vld_25_17 = out_chan_dep_vld_vec_25[16];
    assign dep_chan_data_25_17 = out_chan_dep_data_25;
    assign token_25_17 = token_out_vec_25[16];
    assign dep_chan_vld_25_18 = out_chan_dep_vld_vec_25[17];
    assign dep_chan_data_25_18 = out_chan_dep_data_25;
    assign token_25_18 = token_out_vec_25[17];
    assign dep_chan_vld_25_19 = out_chan_dep_vld_vec_25[18];
    assign dep_chan_data_25_19 = out_chan_dep_data_25;
    assign token_25_19 = token_out_vec_25[18];
    assign dep_chan_vld_25_20 = out_chan_dep_vld_vec_25[19];
    assign dep_chan_data_25_20 = out_chan_dep_data_25;
    assign token_25_20 = token_out_vec_25[19];
    assign dep_chan_vld_25_21 = out_chan_dep_vld_vec_25[20];
    assign dep_chan_data_25_21 = out_chan_dep_data_25;
    assign token_25_21 = token_out_vec_25[20];
    assign dep_chan_vld_25_22 = out_chan_dep_vld_vec_25[21];
    assign dep_chan_data_25_22 = out_chan_dep_data_25;
    assign token_25_22 = token_out_vec_25[21];
    assign dep_chan_vld_25_23 = out_chan_dep_vld_vec_25[22];
    assign dep_chan_data_25_23 = out_chan_dep_data_25;
    assign token_25_23 = token_out_vec_25[22];
    assign dep_chan_vld_25_27 = out_chan_dep_vld_vec_25[23];
    assign dep_chan_data_25_27 = out_chan_dep_data_25;
    assign token_25_27 = token_out_vec_25[23];
    assign dep_chan_vld_25_28 = out_chan_dep_vld_vec_25[24];
    assign dep_chan_data_25_28 = out_chan_dep_data_25;
    assign token_25_28 = token_out_vec_25[24];
    assign dep_chan_vld_25_29 = out_chan_dep_vld_vec_25[25];
    assign dep_chan_data_25_29 = out_chan_dep_data_25;
    assign token_25_29 = token_out_vec_25[25];
    assign dep_chan_vld_25_30 = out_chan_dep_vld_vec_25[26];
    assign dep_chan_data_25_30 = out_chan_dep_data_25;
    assign token_25_30 = token_out_vec_25[26];
    assign dep_chan_vld_25_31 = out_chan_dep_vld_vec_25[27];
    assign dep_chan_data_25_31 = out_chan_dep_data_25;
    assign token_25_31 = token_out_vec_25[27];
    assign dep_chan_vld_25_32 = out_chan_dep_vld_vec_25[28];
    assign dep_chan_data_25_32 = out_chan_dep_data_25;
    assign token_25_32 = token_out_vec_25[28];
    assign dep_chan_vld_25_33 = out_chan_dep_vld_vec_25[29];
    assign dep_chan_data_25_33 = out_chan_dep_data_25;
    assign token_25_33 = token_out_vec_25[29];
    assign dep_chan_vld_25_34 = out_chan_dep_vld_vec_25[30];
    assign dep_chan_data_25_34 = out_chan_dep_data_25;
    assign token_25_34 = token_out_vec_25[30];
    assign dep_chan_vld_25_35 = out_chan_dep_vld_vec_25[31];
    assign dep_chan_data_25_35 = out_chan_dep_data_25;
    assign token_25_35 = token_out_vec_25[31];
    assign dep_chan_vld_25_36 = out_chan_dep_vld_vec_25[32];
    assign dep_chan_data_25_36 = out_chan_dep_data_25;
    assign token_25_36 = token_out_vec_25[32];

    // Process: ProcessingElement_21_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 26, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_26 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_26),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_26),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_26),
        .token_in_vec(token_in_vec_26),
        .dl_detect_in(dl_detect_out),
        .origin(origin[26]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_26),
        .out_chan_dep_data(out_chan_dep_data_26),
        .token_out_vec(token_out_vec_26),
        .dl_detect_out(dl_in_vec[26]));

    assign proc_26_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_20_blk_n) | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_20_blk_n) | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_WriteC_Flattened_fu_179.cPipes_20_blk_n);
    assign proc_26_data_PIPO_blk[0] = 1'b0;
    assign proc_26_start_FIFO_blk[0] = 1'b0;
    assign proc_26_TLF_FIFO_blk[0] = 1'b0;
    assign proc_26_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_26_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_26[0] = dl_detect_out ? proc_dep_vld_vec_26_reg[0] : (proc_26_data_FIFO_blk[0] | proc_26_data_PIPO_blk[0] | proc_26_start_FIFO_blk[0] | proc_26_TLF_FIFO_blk[0] | proc_26_input_sync_blk[0] | proc_26_output_sync_blk[0]);
    assign proc_26_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_21_blk_n) | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_21_blk_n) | (~ProcessingElement_21_U0.grp_ProcessingElement_21_Pipeline_WriteC_Flattened_fu_179.cPipes_21_blk_n);
    assign proc_26_data_PIPO_blk[1] = 1'b0;
    assign proc_26_start_FIFO_blk[1] = 1'b0;
    assign proc_26_TLF_FIFO_blk[1] = 1'b0;
    assign proc_26_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_26_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_26[1] = dl_detect_out ? proc_dep_vld_vec_26_reg[1] : (proc_26_data_FIFO_blk[1] | proc_26_data_PIPO_blk[1] | proc_26_start_FIFO_blk[1] | proc_26_TLF_FIFO_blk[1] | proc_26_input_sync_blk[1] | proc_26_output_sync_blk[1]);
    assign proc_26_data_FIFO_blk[2] = 1'b0;
    assign proc_26_data_PIPO_blk[2] = 1'b0;
    assign proc_26_start_FIFO_blk[2] = 1'b0;
    assign proc_26_TLF_FIFO_blk[2] = 1'b0;
    assign proc_26_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_26_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_26[2] = dl_detect_out ? proc_dep_vld_vec_26_reg[2] : (proc_26_data_FIFO_blk[2] | proc_26_data_PIPO_blk[2] | proc_26_start_FIFO_blk[2] | proc_26_TLF_FIFO_blk[2] | proc_26_input_sync_blk[2] | proc_26_output_sync_blk[2]);
    assign proc_26_data_FIFO_blk[3] = 1'b0;
    assign proc_26_data_PIPO_blk[3] = 1'b0;
    assign proc_26_start_FIFO_blk[3] = 1'b0;
    assign proc_26_TLF_FIFO_blk[3] = 1'b0;
    assign proc_26_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_26_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_26[3] = dl_detect_out ? proc_dep_vld_vec_26_reg[3] : (proc_26_data_FIFO_blk[3] | proc_26_data_PIPO_blk[3] | proc_26_start_FIFO_blk[3] | proc_26_TLF_FIFO_blk[3] | proc_26_input_sync_blk[3] | proc_26_output_sync_blk[3]);
    assign proc_26_data_FIFO_blk[4] = 1'b0;
    assign proc_26_data_PIPO_blk[4] = 1'b0;
    assign proc_26_start_FIFO_blk[4] = 1'b0;
    assign proc_26_TLF_FIFO_blk[4] = 1'b0;
    assign proc_26_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_26_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_26[4] = dl_detect_out ? proc_dep_vld_vec_26_reg[4] : (proc_26_data_FIFO_blk[4] | proc_26_data_PIPO_blk[4] | proc_26_start_FIFO_blk[4] | proc_26_TLF_FIFO_blk[4] | proc_26_input_sync_blk[4] | proc_26_output_sync_blk[4]);
    assign proc_26_data_FIFO_blk[5] = 1'b0;
    assign proc_26_data_PIPO_blk[5] = 1'b0;
    assign proc_26_start_FIFO_blk[5] = 1'b0;
    assign proc_26_TLF_FIFO_blk[5] = 1'b0;
    assign proc_26_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_26_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_26[5] = dl_detect_out ? proc_dep_vld_vec_26_reg[5] : (proc_26_data_FIFO_blk[5] | proc_26_data_PIPO_blk[5] | proc_26_start_FIFO_blk[5] | proc_26_TLF_FIFO_blk[5] | proc_26_input_sync_blk[5] | proc_26_output_sync_blk[5]);
    assign proc_26_data_FIFO_blk[6] = 1'b0;
    assign proc_26_data_PIPO_blk[6] = 1'b0;
    assign proc_26_start_FIFO_blk[6] = 1'b0;
    assign proc_26_TLF_FIFO_blk[6] = 1'b0;
    assign proc_26_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_26_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_26[6] = dl_detect_out ? proc_dep_vld_vec_26_reg[6] : (proc_26_data_FIFO_blk[6] | proc_26_data_PIPO_blk[6] | proc_26_start_FIFO_blk[6] | proc_26_TLF_FIFO_blk[6] | proc_26_input_sync_blk[6] | proc_26_output_sync_blk[6]);
    assign proc_26_data_FIFO_blk[7] = 1'b0;
    assign proc_26_data_PIPO_blk[7] = 1'b0;
    assign proc_26_start_FIFO_blk[7] = 1'b0;
    assign proc_26_TLF_FIFO_blk[7] = 1'b0;
    assign proc_26_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_26_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_26[7] = dl_detect_out ? proc_dep_vld_vec_26_reg[7] : (proc_26_data_FIFO_blk[7] | proc_26_data_PIPO_blk[7] | proc_26_start_FIFO_blk[7] | proc_26_TLF_FIFO_blk[7] | proc_26_input_sync_blk[7] | proc_26_output_sync_blk[7]);
    assign proc_26_data_FIFO_blk[8] = 1'b0;
    assign proc_26_data_PIPO_blk[8] = 1'b0;
    assign proc_26_start_FIFO_blk[8] = 1'b0;
    assign proc_26_TLF_FIFO_blk[8] = 1'b0;
    assign proc_26_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_26_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_26[8] = dl_detect_out ? proc_dep_vld_vec_26_reg[8] : (proc_26_data_FIFO_blk[8] | proc_26_data_PIPO_blk[8] | proc_26_start_FIFO_blk[8] | proc_26_TLF_FIFO_blk[8] | proc_26_input_sync_blk[8] | proc_26_output_sync_blk[8]);
    assign proc_26_data_FIFO_blk[9] = 1'b0;
    assign proc_26_data_PIPO_blk[9] = 1'b0;
    assign proc_26_start_FIFO_blk[9] = 1'b0;
    assign proc_26_TLF_FIFO_blk[9] = 1'b0;
    assign proc_26_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_26_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_26[9] = dl_detect_out ? proc_dep_vld_vec_26_reg[9] : (proc_26_data_FIFO_blk[9] | proc_26_data_PIPO_blk[9] | proc_26_start_FIFO_blk[9] | proc_26_TLF_FIFO_blk[9] | proc_26_input_sync_blk[9] | proc_26_output_sync_blk[9]);
    assign proc_26_data_FIFO_blk[10] = 1'b0;
    assign proc_26_data_PIPO_blk[10] = 1'b0;
    assign proc_26_start_FIFO_blk[10] = 1'b0;
    assign proc_26_TLF_FIFO_blk[10] = 1'b0;
    assign proc_26_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_26_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_26[10] = dl_detect_out ? proc_dep_vld_vec_26_reg[10] : (proc_26_data_FIFO_blk[10] | proc_26_data_PIPO_blk[10] | proc_26_start_FIFO_blk[10] | proc_26_TLF_FIFO_blk[10] | proc_26_input_sync_blk[10] | proc_26_output_sync_blk[10]);
    assign proc_26_data_FIFO_blk[11] = 1'b0;
    assign proc_26_data_PIPO_blk[11] = 1'b0;
    assign proc_26_start_FIFO_blk[11] = 1'b0;
    assign proc_26_TLF_FIFO_blk[11] = 1'b0;
    assign proc_26_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_26_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_26[11] = dl_detect_out ? proc_dep_vld_vec_26_reg[11] : (proc_26_data_FIFO_blk[11] | proc_26_data_PIPO_blk[11] | proc_26_start_FIFO_blk[11] | proc_26_TLF_FIFO_blk[11] | proc_26_input_sync_blk[11] | proc_26_output_sync_blk[11]);
    assign proc_26_data_FIFO_blk[12] = 1'b0;
    assign proc_26_data_PIPO_blk[12] = 1'b0;
    assign proc_26_start_FIFO_blk[12] = 1'b0;
    assign proc_26_TLF_FIFO_blk[12] = 1'b0;
    assign proc_26_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_26_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_26[12] = dl_detect_out ? proc_dep_vld_vec_26_reg[12] : (proc_26_data_FIFO_blk[12] | proc_26_data_PIPO_blk[12] | proc_26_start_FIFO_blk[12] | proc_26_TLF_FIFO_blk[12] | proc_26_input_sync_blk[12] | proc_26_output_sync_blk[12]);
    assign proc_26_data_FIFO_blk[13] = 1'b0;
    assign proc_26_data_PIPO_blk[13] = 1'b0;
    assign proc_26_start_FIFO_blk[13] = 1'b0;
    assign proc_26_TLF_FIFO_blk[13] = 1'b0;
    assign proc_26_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_26_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_26[13] = dl_detect_out ? proc_dep_vld_vec_26_reg[13] : (proc_26_data_FIFO_blk[13] | proc_26_data_PIPO_blk[13] | proc_26_start_FIFO_blk[13] | proc_26_TLF_FIFO_blk[13] | proc_26_input_sync_blk[13] | proc_26_output_sync_blk[13]);
    assign proc_26_data_FIFO_blk[14] = 1'b0;
    assign proc_26_data_PIPO_blk[14] = 1'b0;
    assign proc_26_start_FIFO_blk[14] = 1'b0;
    assign proc_26_TLF_FIFO_blk[14] = 1'b0;
    assign proc_26_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_26_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_26[14] = dl_detect_out ? proc_dep_vld_vec_26_reg[14] : (proc_26_data_FIFO_blk[14] | proc_26_data_PIPO_blk[14] | proc_26_start_FIFO_blk[14] | proc_26_TLF_FIFO_blk[14] | proc_26_input_sync_blk[14] | proc_26_output_sync_blk[14]);
    assign proc_26_data_FIFO_blk[15] = 1'b0;
    assign proc_26_data_PIPO_blk[15] = 1'b0;
    assign proc_26_start_FIFO_blk[15] = 1'b0;
    assign proc_26_TLF_FIFO_blk[15] = 1'b0;
    assign proc_26_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_26_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_26[15] = dl_detect_out ? proc_dep_vld_vec_26_reg[15] : (proc_26_data_FIFO_blk[15] | proc_26_data_PIPO_blk[15] | proc_26_start_FIFO_blk[15] | proc_26_TLF_FIFO_blk[15] | proc_26_input_sync_blk[15] | proc_26_output_sync_blk[15]);
    assign proc_26_data_FIFO_blk[16] = 1'b0;
    assign proc_26_data_PIPO_blk[16] = 1'b0;
    assign proc_26_start_FIFO_blk[16] = 1'b0;
    assign proc_26_TLF_FIFO_blk[16] = 1'b0;
    assign proc_26_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_26_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_26[16] = dl_detect_out ? proc_dep_vld_vec_26_reg[16] : (proc_26_data_FIFO_blk[16] | proc_26_data_PIPO_blk[16] | proc_26_start_FIFO_blk[16] | proc_26_TLF_FIFO_blk[16] | proc_26_input_sync_blk[16] | proc_26_output_sync_blk[16]);
    assign proc_26_data_FIFO_blk[17] = 1'b0;
    assign proc_26_data_PIPO_blk[17] = 1'b0;
    assign proc_26_start_FIFO_blk[17] = 1'b0;
    assign proc_26_TLF_FIFO_blk[17] = 1'b0;
    assign proc_26_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_26_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_26[17] = dl_detect_out ? proc_dep_vld_vec_26_reg[17] : (proc_26_data_FIFO_blk[17] | proc_26_data_PIPO_blk[17] | proc_26_start_FIFO_blk[17] | proc_26_TLF_FIFO_blk[17] | proc_26_input_sync_blk[17] | proc_26_output_sync_blk[17]);
    assign proc_26_data_FIFO_blk[18] = 1'b0;
    assign proc_26_data_PIPO_blk[18] = 1'b0;
    assign proc_26_start_FIFO_blk[18] = 1'b0;
    assign proc_26_TLF_FIFO_blk[18] = 1'b0;
    assign proc_26_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_26_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_26[18] = dl_detect_out ? proc_dep_vld_vec_26_reg[18] : (proc_26_data_FIFO_blk[18] | proc_26_data_PIPO_blk[18] | proc_26_start_FIFO_blk[18] | proc_26_TLF_FIFO_blk[18] | proc_26_input_sync_blk[18] | proc_26_output_sync_blk[18]);
    assign proc_26_data_FIFO_blk[19] = 1'b0;
    assign proc_26_data_PIPO_blk[19] = 1'b0;
    assign proc_26_start_FIFO_blk[19] = 1'b0;
    assign proc_26_TLF_FIFO_blk[19] = 1'b0;
    assign proc_26_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_26_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_26[19] = dl_detect_out ? proc_dep_vld_vec_26_reg[19] : (proc_26_data_FIFO_blk[19] | proc_26_data_PIPO_blk[19] | proc_26_start_FIFO_blk[19] | proc_26_TLF_FIFO_blk[19] | proc_26_input_sync_blk[19] | proc_26_output_sync_blk[19]);
    assign proc_26_data_FIFO_blk[20] = 1'b0;
    assign proc_26_data_PIPO_blk[20] = 1'b0;
    assign proc_26_start_FIFO_blk[20] = 1'b0;
    assign proc_26_TLF_FIFO_blk[20] = 1'b0;
    assign proc_26_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_26_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_26[20] = dl_detect_out ? proc_dep_vld_vec_26_reg[20] : (proc_26_data_FIFO_blk[20] | proc_26_data_PIPO_blk[20] | proc_26_start_FIFO_blk[20] | proc_26_TLF_FIFO_blk[20] | proc_26_input_sync_blk[20] | proc_26_output_sync_blk[20]);
    assign proc_26_data_FIFO_blk[21] = 1'b0;
    assign proc_26_data_PIPO_blk[21] = 1'b0;
    assign proc_26_start_FIFO_blk[21] = 1'b0;
    assign proc_26_TLF_FIFO_blk[21] = 1'b0;
    assign proc_26_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_26_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_26[21] = dl_detect_out ? proc_dep_vld_vec_26_reg[21] : (proc_26_data_FIFO_blk[21] | proc_26_data_PIPO_blk[21] | proc_26_start_FIFO_blk[21] | proc_26_TLF_FIFO_blk[21] | proc_26_input_sync_blk[21] | proc_26_output_sync_blk[21]);
    assign proc_26_data_FIFO_blk[22] = 1'b0;
    assign proc_26_data_PIPO_blk[22] = 1'b0;
    assign proc_26_start_FIFO_blk[22] = 1'b0;
    assign proc_26_TLF_FIFO_blk[22] = 1'b0;
    assign proc_26_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_26_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_26[22] = dl_detect_out ? proc_dep_vld_vec_26_reg[22] : (proc_26_data_FIFO_blk[22] | proc_26_data_PIPO_blk[22] | proc_26_start_FIFO_blk[22] | proc_26_TLF_FIFO_blk[22] | proc_26_input_sync_blk[22] | proc_26_output_sync_blk[22]);
    assign proc_26_data_FIFO_blk[23] = 1'b0;
    assign proc_26_data_PIPO_blk[23] = 1'b0;
    assign proc_26_start_FIFO_blk[23] = 1'b0;
    assign proc_26_TLF_FIFO_blk[23] = 1'b0;
    assign proc_26_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_26_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_26[23] = dl_detect_out ? proc_dep_vld_vec_26_reg[23] : (proc_26_data_FIFO_blk[23] | proc_26_data_PIPO_blk[23] | proc_26_start_FIFO_blk[23] | proc_26_TLF_FIFO_blk[23] | proc_26_input_sync_blk[23] | proc_26_output_sync_blk[23]);
    assign proc_26_data_FIFO_blk[24] = 1'b0;
    assign proc_26_data_PIPO_blk[24] = 1'b0;
    assign proc_26_start_FIFO_blk[24] = 1'b0;
    assign proc_26_TLF_FIFO_blk[24] = 1'b0;
    assign proc_26_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_26_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_26[24] = dl_detect_out ? proc_dep_vld_vec_26_reg[24] : (proc_26_data_FIFO_blk[24] | proc_26_data_PIPO_blk[24] | proc_26_start_FIFO_blk[24] | proc_26_TLF_FIFO_blk[24] | proc_26_input_sync_blk[24] | proc_26_output_sync_blk[24]);
    assign proc_26_data_FIFO_blk[25] = 1'b0;
    assign proc_26_data_PIPO_blk[25] = 1'b0;
    assign proc_26_start_FIFO_blk[25] = 1'b0;
    assign proc_26_TLF_FIFO_blk[25] = 1'b0;
    assign proc_26_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_26_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_26[25] = dl_detect_out ? proc_dep_vld_vec_26_reg[25] : (proc_26_data_FIFO_blk[25] | proc_26_data_PIPO_blk[25] | proc_26_start_FIFO_blk[25] | proc_26_TLF_FIFO_blk[25] | proc_26_input_sync_blk[25] | proc_26_output_sync_blk[25]);
    assign proc_26_data_FIFO_blk[26] = 1'b0;
    assign proc_26_data_PIPO_blk[26] = 1'b0;
    assign proc_26_start_FIFO_blk[26] = 1'b0;
    assign proc_26_TLF_FIFO_blk[26] = 1'b0;
    assign proc_26_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_26_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_26[26] = dl_detect_out ? proc_dep_vld_vec_26_reg[26] : (proc_26_data_FIFO_blk[26] | proc_26_data_PIPO_blk[26] | proc_26_start_FIFO_blk[26] | proc_26_TLF_FIFO_blk[26] | proc_26_input_sync_blk[26] | proc_26_output_sync_blk[26]);
    assign proc_26_data_FIFO_blk[27] = 1'b0;
    assign proc_26_data_PIPO_blk[27] = 1'b0;
    assign proc_26_start_FIFO_blk[27] = 1'b0;
    assign proc_26_TLF_FIFO_blk[27] = 1'b0;
    assign proc_26_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_26_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_26[27] = dl_detect_out ? proc_dep_vld_vec_26_reg[27] : (proc_26_data_FIFO_blk[27] | proc_26_data_PIPO_blk[27] | proc_26_start_FIFO_blk[27] | proc_26_TLF_FIFO_blk[27] | proc_26_input_sync_blk[27] | proc_26_output_sync_blk[27]);
    assign proc_26_data_FIFO_blk[28] = 1'b0;
    assign proc_26_data_PIPO_blk[28] = 1'b0;
    assign proc_26_start_FIFO_blk[28] = 1'b0;
    assign proc_26_TLF_FIFO_blk[28] = 1'b0;
    assign proc_26_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_26_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_26[28] = dl_detect_out ? proc_dep_vld_vec_26_reg[28] : (proc_26_data_FIFO_blk[28] | proc_26_data_PIPO_blk[28] | proc_26_start_FIFO_blk[28] | proc_26_TLF_FIFO_blk[28] | proc_26_input_sync_blk[28] | proc_26_output_sync_blk[28]);
    assign proc_26_data_FIFO_blk[29] = 1'b0;
    assign proc_26_data_PIPO_blk[29] = 1'b0;
    assign proc_26_start_FIFO_blk[29] = 1'b0;
    assign proc_26_TLF_FIFO_blk[29] = 1'b0;
    assign proc_26_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_26_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_26[29] = dl_detect_out ? proc_dep_vld_vec_26_reg[29] : (proc_26_data_FIFO_blk[29] | proc_26_data_PIPO_blk[29] | proc_26_start_FIFO_blk[29] | proc_26_TLF_FIFO_blk[29] | proc_26_input_sync_blk[29] | proc_26_output_sync_blk[29]);
    assign proc_26_data_FIFO_blk[30] = 1'b0;
    assign proc_26_data_PIPO_blk[30] = 1'b0;
    assign proc_26_start_FIFO_blk[30] = 1'b0;
    assign proc_26_TLF_FIFO_blk[30] = 1'b0;
    assign proc_26_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_26_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_26[30] = dl_detect_out ? proc_dep_vld_vec_26_reg[30] : (proc_26_data_FIFO_blk[30] | proc_26_data_PIPO_blk[30] | proc_26_start_FIFO_blk[30] | proc_26_TLF_FIFO_blk[30] | proc_26_input_sync_blk[30] | proc_26_output_sync_blk[30]);
    assign proc_26_data_FIFO_blk[31] = 1'b0;
    assign proc_26_data_PIPO_blk[31] = 1'b0;
    assign proc_26_start_FIFO_blk[31] = 1'b0;
    assign proc_26_TLF_FIFO_blk[31] = 1'b0;
    assign proc_26_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_26_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_26[31] = dl_detect_out ? proc_dep_vld_vec_26_reg[31] : (proc_26_data_FIFO_blk[31] | proc_26_data_PIPO_blk[31] | proc_26_start_FIFO_blk[31] | proc_26_TLF_FIFO_blk[31] | proc_26_input_sync_blk[31] | proc_26_output_sync_blk[31]);
    assign proc_26_data_FIFO_blk[32] = 1'b0;
    assign proc_26_data_PIPO_blk[32] = 1'b0;
    assign proc_26_start_FIFO_blk[32] = 1'b0;
    assign proc_26_TLF_FIFO_blk[32] = 1'b0;
    assign proc_26_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_21_U0_ap_ready & ProcessingElement_21_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_26_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_26[32] = dl_detect_out ? proc_dep_vld_vec_26_reg[32] : (proc_26_data_FIFO_blk[32] | proc_26_data_PIPO_blk[32] | proc_26_start_FIFO_blk[32] | proc_26_TLF_FIFO_blk[32] | proc_26_input_sync_blk[32] | proc_26_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_26_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_26_reg <= proc_dep_vld_vec_26;
        end
    end
    assign in_chan_dep_vld_vec_26[0] = dep_chan_vld_0_26;
    assign in_chan_dep_data_vec_26[39 : 0] = dep_chan_data_0_26;
    assign token_in_vec_26[0] = token_0_26;
    assign in_chan_dep_vld_vec_26[1] = dep_chan_vld_1_26;
    assign in_chan_dep_data_vec_26[79 : 40] = dep_chan_data_1_26;
    assign token_in_vec_26[1] = token_1_26;
    assign in_chan_dep_vld_vec_26[2] = dep_chan_vld_3_26;
    assign in_chan_dep_data_vec_26[119 : 80] = dep_chan_data_3_26;
    assign token_in_vec_26[2] = token_3_26;
    assign in_chan_dep_vld_vec_26[3] = dep_chan_vld_6_26;
    assign in_chan_dep_data_vec_26[159 : 120] = dep_chan_data_6_26;
    assign token_in_vec_26[3] = token_6_26;
    assign in_chan_dep_vld_vec_26[4] = dep_chan_vld_7_26;
    assign in_chan_dep_data_vec_26[199 : 160] = dep_chan_data_7_26;
    assign token_in_vec_26[4] = token_7_26;
    assign in_chan_dep_vld_vec_26[5] = dep_chan_vld_8_26;
    assign in_chan_dep_data_vec_26[239 : 200] = dep_chan_data_8_26;
    assign token_in_vec_26[5] = token_8_26;
    assign in_chan_dep_vld_vec_26[6] = dep_chan_vld_9_26;
    assign in_chan_dep_data_vec_26[279 : 240] = dep_chan_data_9_26;
    assign token_in_vec_26[6] = token_9_26;
    assign in_chan_dep_vld_vec_26[7] = dep_chan_vld_10_26;
    assign in_chan_dep_data_vec_26[319 : 280] = dep_chan_data_10_26;
    assign token_in_vec_26[7] = token_10_26;
    assign in_chan_dep_vld_vec_26[8] = dep_chan_vld_11_26;
    assign in_chan_dep_data_vec_26[359 : 320] = dep_chan_data_11_26;
    assign token_in_vec_26[8] = token_11_26;
    assign in_chan_dep_vld_vec_26[9] = dep_chan_vld_12_26;
    assign in_chan_dep_data_vec_26[399 : 360] = dep_chan_data_12_26;
    assign token_in_vec_26[9] = token_12_26;
    assign in_chan_dep_vld_vec_26[10] = dep_chan_vld_13_26;
    assign in_chan_dep_data_vec_26[439 : 400] = dep_chan_data_13_26;
    assign token_in_vec_26[10] = token_13_26;
    assign in_chan_dep_vld_vec_26[11] = dep_chan_vld_14_26;
    assign in_chan_dep_data_vec_26[479 : 440] = dep_chan_data_14_26;
    assign token_in_vec_26[11] = token_14_26;
    assign in_chan_dep_vld_vec_26[12] = dep_chan_vld_15_26;
    assign in_chan_dep_data_vec_26[519 : 480] = dep_chan_data_15_26;
    assign token_in_vec_26[12] = token_15_26;
    assign in_chan_dep_vld_vec_26[13] = dep_chan_vld_16_26;
    assign in_chan_dep_data_vec_26[559 : 520] = dep_chan_data_16_26;
    assign token_in_vec_26[13] = token_16_26;
    assign in_chan_dep_vld_vec_26[14] = dep_chan_vld_17_26;
    assign in_chan_dep_data_vec_26[599 : 560] = dep_chan_data_17_26;
    assign token_in_vec_26[14] = token_17_26;
    assign in_chan_dep_vld_vec_26[15] = dep_chan_vld_18_26;
    assign in_chan_dep_data_vec_26[639 : 600] = dep_chan_data_18_26;
    assign token_in_vec_26[15] = token_18_26;
    assign in_chan_dep_vld_vec_26[16] = dep_chan_vld_19_26;
    assign in_chan_dep_data_vec_26[679 : 640] = dep_chan_data_19_26;
    assign token_in_vec_26[16] = token_19_26;
    assign in_chan_dep_vld_vec_26[17] = dep_chan_vld_20_26;
    assign in_chan_dep_data_vec_26[719 : 680] = dep_chan_data_20_26;
    assign token_in_vec_26[17] = token_20_26;
    assign in_chan_dep_vld_vec_26[18] = dep_chan_vld_21_26;
    assign in_chan_dep_data_vec_26[759 : 720] = dep_chan_data_21_26;
    assign token_in_vec_26[18] = token_21_26;
    assign in_chan_dep_vld_vec_26[19] = dep_chan_vld_22_26;
    assign in_chan_dep_data_vec_26[799 : 760] = dep_chan_data_22_26;
    assign token_in_vec_26[19] = token_22_26;
    assign in_chan_dep_vld_vec_26[20] = dep_chan_vld_23_26;
    assign in_chan_dep_data_vec_26[839 : 800] = dep_chan_data_23_26;
    assign token_in_vec_26[20] = token_23_26;
    assign in_chan_dep_vld_vec_26[21] = dep_chan_vld_24_26;
    assign in_chan_dep_data_vec_26[879 : 840] = dep_chan_data_24_26;
    assign token_in_vec_26[21] = token_24_26;
    assign in_chan_dep_vld_vec_26[22] = dep_chan_vld_25_26;
    assign in_chan_dep_data_vec_26[919 : 880] = dep_chan_data_25_26;
    assign token_in_vec_26[22] = token_25_26;
    assign in_chan_dep_vld_vec_26[23] = dep_chan_vld_27_26;
    assign in_chan_dep_data_vec_26[959 : 920] = dep_chan_data_27_26;
    assign token_in_vec_26[23] = token_27_26;
    assign in_chan_dep_vld_vec_26[24] = dep_chan_vld_28_26;
    assign in_chan_dep_data_vec_26[999 : 960] = dep_chan_data_28_26;
    assign token_in_vec_26[24] = token_28_26;
    assign in_chan_dep_vld_vec_26[25] = dep_chan_vld_29_26;
    assign in_chan_dep_data_vec_26[1039 : 1000] = dep_chan_data_29_26;
    assign token_in_vec_26[25] = token_29_26;
    assign in_chan_dep_vld_vec_26[26] = dep_chan_vld_30_26;
    assign in_chan_dep_data_vec_26[1079 : 1040] = dep_chan_data_30_26;
    assign token_in_vec_26[26] = token_30_26;
    assign in_chan_dep_vld_vec_26[27] = dep_chan_vld_31_26;
    assign in_chan_dep_data_vec_26[1119 : 1080] = dep_chan_data_31_26;
    assign token_in_vec_26[27] = token_31_26;
    assign in_chan_dep_vld_vec_26[28] = dep_chan_vld_32_26;
    assign in_chan_dep_data_vec_26[1159 : 1120] = dep_chan_data_32_26;
    assign token_in_vec_26[28] = token_32_26;
    assign in_chan_dep_vld_vec_26[29] = dep_chan_vld_33_26;
    assign in_chan_dep_data_vec_26[1199 : 1160] = dep_chan_data_33_26;
    assign token_in_vec_26[29] = token_33_26;
    assign in_chan_dep_vld_vec_26[30] = dep_chan_vld_34_26;
    assign in_chan_dep_data_vec_26[1239 : 1200] = dep_chan_data_34_26;
    assign token_in_vec_26[30] = token_34_26;
    assign in_chan_dep_vld_vec_26[31] = dep_chan_vld_35_26;
    assign in_chan_dep_data_vec_26[1279 : 1240] = dep_chan_data_35_26;
    assign token_in_vec_26[31] = token_35_26;
    assign in_chan_dep_vld_vec_26[32] = dep_chan_vld_36_26;
    assign in_chan_dep_data_vec_26[1319 : 1280] = dep_chan_data_36_26;
    assign token_in_vec_26[32] = token_36_26;
    assign dep_chan_vld_26_25 = out_chan_dep_vld_vec_26[0];
    assign dep_chan_data_26_25 = out_chan_dep_data_26;
    assign token_26_25 = token_out_vec_26[0];
    assign dep_chan_vld_26_27 = out_chan_dep_vld_vec_26[1];
    assign dep_chan_data_26_27 = out_chan_dep_data_26;
    assign token_26_27 = token_out_vec_26[1];
    assign dep_chan_vld_26_0 = out_chan_dep_vld_vec_26[2];
    assign dep_chan_data_26_0 = out_chan_dep_data_26;
    assign token_26_0 = token_out_vec_26[2];
    assign dep_chan_vld_26_1 = out_chan_dep_vld_vec_26[3];
    assign dep_chan_data_26_1 = out_chan_dep_data_26;
    assign token_26_1 = token_out_vec_26[3];
    assign dep_chan_vld_26_3 = out_chan_dep_vld_vec_26[4];
    assign dep_chan_data_26_3 = out_chan_dep_data_26;
    assign token_26_3 = token_out_vec_26[4];
    assign dep_chan_vld_26_6 = out_chan_dep_vld_vec_26[5];
    assign dep_chan_data_26_6 = out_chan_dep_data_26;
    assign token_26_6 = token_out_vec_26[5];
    assign dep_chan_vld_26_7 = out_chan_dep_vld_vec_26[6];
    assign dep_chan_data_26_7 = out_chan_dep_data_26;
    assign token_26_7 = token_out_vec_26[6];
    assign dep_chan_vld_26_8 = out_chan_dep_vld_vec_26[7];
    assign dep_chan_data_26_8 = out_chan_dep_data_26;
    assign token_26_8 = token_out_vec_26[7];
    assign dep_chan_vld_26_9 = out_chan_dep_vld_vec_26[8];
    assign dep_chan_data_26_9 = out_chan_dep_data_26;
    assign token_26_9 = token_out_vec_26[8];
    assign dep_chan_vld_26_10 = out_chan_dep_vld_vec_26[9];
    assign dep_chan_data_26_10 = out_chan_dep_data_26;
    assign token_26_10 = token_out_vec_26[9];
    assign dep_chan_vld_26_11 = out_chan_dep_vld_vec_26[10];
    assign dep_chan_data_26_11 = out_chan_dep_data_26;
    assign token_26_11 = token_out_vec_26[10];
    assign dep_chan_vld_26_12 = out_chan_dep_vld_vec_26[11];
    assign dep_chan_data_26_12 = out_chan_dep_data_26;
    assign token_26_12 = token_out_vec_26[11];
    assign dep_chan_vld_26_13 = out_chan_dep_vld_vec_26[12];
    assign dep_chan_data_26_13 = out_chan_dep_data_26;
    assign token_26_13 = token_out_vec_26[12];
    assign dep_chan_vld_26_14 = out_chan_dep_vld_vec_26[13];
    assign dep_chan_data_26_14 = out_chan_dep_data_26;
    assign token_26_14 = token_out_vec_26[13];
    assign dep_chan_vld_26_15 = out_chan_dep_vld_vec_26[14];
    assign dep_chan_data_26_15 = out_chan_dep_data_26;
    assign token_26_15 = token_out_vec_26[14];
    assign dep_chan_vld_26_16 = out_chan_dep_vld_vec_26[15];
    assign dep_chan_data_26_16 = out_chan_dep_data_26;
    assign token_26_16 = token_out_vec_26[15];
    assign dep_chan_vld_26_17 = out_chan_dep_vld_vec_26[16];
    assign dep_chan_data_26_17 = out_chan_dep_data_26;
    assign token_26_17 = token_out_vec_26[16];
    assign dep_chan_vld_26_18 = out_chan_dep_vld_vec_26[17];
    assign dep_chan_data_26_18 = out_chan_dep_data_26;
    assign token_26_18 = token_out_vec_26[17];
    assign dep_chan_vld_26_19 = out_chan_dep_vld_vec_26[18];
    assign dep_chan_data_26_19 = out_chan_dep_data_26;
    assign token_26_19 = token_out_vec_26[18];
    assign dep_chan_vld_26_20 = out_chan_dep_vld_vec_26[19];
    assign dep_chan_data_26_20 = out_chan_dep_data_26;
    assign token_26_20 = token_out_vec_26[19];
    assign dep_chan_vld_26_21 = out_chan_dep_vld_vec_26[20];
    assign dep_chan_data_26_21 = out_chan_dep_data_26;
    assign token_26_21 = token_out_vec_26[20];
    assign dep_chan_vld_26_22 = out_chan_dep_vld_vec_26[21];
    assign dep_chan_data_26_22 = out_chan_dep_data_26;
    assign token_26_22 = token_out_vec_26[21];
    assign dep_chan_vld_26_23 = out_chan_dep_vld_vec_26[22];
    assign dep_chan_data_26_23 = out_chan_dep_data_26;
    assign token_26_23 = token_out_vec_26[22];
    assign dep_chan_vld_26_24 = out_chan_dep_vld_vec_26[23];
    assign dep_chan_data_26_24 = out_chan_dep_data_26;
    assign token_26_24 = token_out_vec_26[23];
    assign dep_chan_vld_26_28 = out_chan_dep_vld_vec_26[24];
    assign dep_chan_data_26_28 = out_chan_dep_data_26;
    assign token_26_28 = token_out_vec_26[24];
    assign dep_chan_vld_26_29 = out_chan_dep_vld_vec_26[25];
    assign dep_chan_data_26_29 = out_chan_dep_data_26;
    assign token_26_29 = token_out_vec_26[25];
    assign dep_chan_vld_26_30 = out_chan_dep_vld_vec_26[26];
    assign dep_chan_data_26_30 = out_chan_dep_data_26;
    assign token_26_30 = token_out_vec_26[26];
    assign dep_chan_vld_26_31 = out_chan_dep_vld_vec_26[27];
    assign dep_chan_data_26_31 = out_chan_dep_data_26;
    assign token_26_31 = token_out_vec_26[27];
    assign dep_chan_vld_26_32 = out_chan_dep_vld_vec_26[28];
    assign dep_chan_data_26_32 = out_chan_dep_data_26;
    assign token_26_32 = token_out_vec_26[28];
    assign dep_chan_vld_26_33 = out_chan_dep_vld_vec_26[29];
    assign dep_chan_data_26_33 = out_chan_dep_data_26;
    assign token_26_33 = token_out_vec_26[29];
    assign dep_chan_vld_26_34 = out_chan_dep_vld_vec_26[30];
    assign dep_chan_data_26_34 = out_chan_dep_data_26;
    assign token_26_34 = token_out_vec_26[30];
    assign dep_chan_vld_26_35 = out_chan_dep_vld_vec_26[31];
    assign dep_chan_data_26_35 = out_chan_dep_data_26;
    assign token_26_35 = token_out_vec_26[31];
    assign dep_chan_vld_26_36 = out_chan_dep_vld_vec_26[32];
    assign dep_chan_data_26_36 = out_chan_dep_data_26;
    assign token_26_36 = token_out_vec_26[32];

    // Process: ProcessingElement_22_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 27, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_27 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_27),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_27),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_27),
        .token_in_vec(token_in_vec_27),
        .dl_detect_in(dl_detect_out),
        .origin(origin[27]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_27),
        .out_chan_dep_data(out_chan_dep_data_27),
        .token_out_vec(token_out_vec_27),
        .dl_detect_out(dl_in_vec[27]));

    assign proc_27_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_21_blk_n) | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_21_blk_n) | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_WriteC_Flattened_fu_179.cPipes_21_blk_n);
    assign proc_27_data_PIPO_blk[0] = 1'b0;
    assign proc_27_start_FIFO_blk[0] = 1'b0;
    assign proc_27_TLF_FIFO_blk[0] = 1'b0;
    assign proc_27_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_27_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_27[0] = dl_detect_out ? proc_dep_vld_vec_27_reg[0] : (proc_27_data_FIFO_blk[0] | proc_27_data_PIPO_blk[0] | proc_27_start_FIFO_blk[0] | proc_27_TLF_FIFO_blk[0] | proc_27_input_sync_blk[0] | proc_27_output_sync_blk[0]);
    assign proc_27_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_22_blk_n) | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_22_blk_n) | (~ProcessingElement_22_U0.grp_ProcessingElement_22_Pipeline_WriteC_Flattened_fu_179.cPipes_22_blk_n);
    assign proc_27_data_PIPO_blk[1] = 1'b0;
    assign proc_27_start_FIFO_blk[1] = 1'b0;
    assign proc_27_TLF_FIFO_blk[1] = 1'b0;
    assign proc_27_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_27_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_27[1] = dl_detect_out ? proc_dep_vld_vec_27_reg[1] : (proc_27_data_FIFO_blk[1] | proc_27_data_PIPO_blk[1] | proc_27_start_FIFO_blk[1] | proc_27_TLF_FIFO_blk[1] | proc_27_input_sync_blk[1] | proc_27_output_sync_blk[1]);
    assign proc_27_data_FIFO_blk[2] = 1'b0;
    assign proc_27_data_PIPO_blk[2] = 1'b0;
    assign proc_27_start_FIFO_blk[2] = 1'b0;
    assign proc_27_TLF_FIFO_blk[2] = 1'b0;
    assign proc_27_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_27_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_27[2] = dl_detect_out ? proc_dep_vld_vec_27_reg[2] : (proc_27_data_FIFO_blk[2] | proc_27_data_PIPO_blk[2] | proc_27_start_FIFO_blk[2] | proc_27_TLF_FIFO_blk[2] | proc_27_input_sync_blk[2] | proc_27_output_sync_blk[2]);
    assign proc_27_data_FIFO_blk[3] = 1'b0;
    assign proc_27_data_PIPO_blk[3] = 1'b0;
    assign proc_27_start_FIFO_blk[3] = 1'b0;
    assign proc_27_TLF_FIFO_blk[3] = 1'b0;
    assign proc_27_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_27_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_27[3] = dl_detect_out ? proc_dep_vld_vec_27_reg[3] : (proc_27_data_FIFO_blk[3] | proc_27_data_PIPO_blk[3] | proc_27_start_FIFO_blk[3] | proc_27_TLF_FIFO_blk[3] | proc_27_input_sync_blk[3] | proc_27_output_sync_blk[3]);
    assign proc_27_data_FIFO_blk[4] = 1'b0;
    assign proc_27_data_PIPO_blk[4] = 1'b0;
    assign proc_27_start_FIFO_blk[4] = 1'b0;
    assign proc_27_TLF_FIFO_blk[4] = 1'b0;
    assign proc_27_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_27_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_27[4] = dl_detect_out ? proc_dep_vld_vec_27_reg[4] : (proc_27_data_FIFO_blk[4] | proc_27_data_PIPO_blk[4] | proc_27_start_FIFO_blk[4] | proc_27_TLF_FIFO_blk[4] | proc_27_input_sync_blk[4] | proc_27_output_sync_blk[4]);
    assign proc_27_data_FIFO_blk[5] = 1'b0;
    assign proc_27_data_PIPO_blk[5] = 1'b0;
    assign proc_27_start_FIFO_blk[5] = 1'b0;
    assign proc_27_TLF_FIFO_blk[5] = 1'b0;
    assign proc_27_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_27_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_27[5] = dl_detect_out ? proc_dep_vld_vec_27_reg[5] : (proc_27_data_FIFO_blk[5] | proc_27_data_PIPO_blk[5] | proc_27_start_FIFO_blk[5] | proc_27_TLF_FIFO_blk[5] | proc_27_input_sync_blk[5] | proc_27_output_sync_blk[5]);
    assign proc_27_data_FIFO_blk[6] = 1'b0;
    assign proc_27_data_PIPO_blk[6] = 1'b0;
    assign proc_27_start_FIFO_blk[6] = 1'b0;
    assign proc_27_TLF_FIFO_blk[6] = 1'b0;
    assign proc_27_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_27_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_27[6] = dl_detect_out ? proc_dep_vld_vec_27_reg[6] : (proc_27_data_FIFO_blk[6] | proc_27_data_PIPO_blk[6] | proc_27_start_FIFO_blk[6] | proc_27_TLF_FIFO_blk[6] | proc_27_input_sync_blk[6] | proc_27_output_sync_blk[6]);
    assign proc_27_data_FIFO_blk[7] = 1'b0;
    assign proc_27_data_PIPO_blk[7] = 1'b0;
    assign proc_27_start_FIFO_blk[7] = 1'b0;
    assign proc_27_TLF_FIFO_blk[7] = 1'b0;
    assign proc_27_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_27_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_27[7] = dl_detect_out ? proc_dep_vld_vec_27_reg[7] : (proc_27_data_FIFO_blk[7] | proc_27_data_PIPO_blk[7] | proc_27_start_FIFO_blk[7] | proc_27_TLF_FIFO_blk[7] | proc_27_input_sync_blk[7] | proc_27_output_sync_blk[7]);
    assign proc_27_data_FIFO_blk[8] = 1'b0;
    assign proc_27_data_PIPO_blk[8] = 1'b0;
    assign proc_27_start_FIFO_blk[8] = 1'b0;
    assign proc_27_TLF_FIFO_blk[8] = 1'b0;
    assign proc_27_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_27_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_27[8] = dl_detect_out ? proc_dep_vld_vec_27_reg[8] : (proc_27_data_FIFO_blk[8] | proc_27_data_PIPO_blk[8] | proc_27_start_FIFO_blk[8] | proc_27_TLF_FIFO_blk[8] | proc_27_input_sync_blk[8] | proc_27_output_sync_blk[8]);
    assign proc_27_data_FIFO_blk[9] = 1'b0;
    assign proc_27_data_PIPO_blk[9] = 1'b0;
    assign proc_27_start_FIFO_blk[9] = 1'b0;
    assign proc_27_TLF_FIFO_blk[9] = 1'b0;
    assign proc_27_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_27_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_27[9] = dl_detect_out ? proc_dep_vld_vec_27_reg[9] : (proc_27_data_FIFO_blk[9] | proc_27_data_PIPO_blk[9] | proc_27_start_FIFO_blk[9] | proc_27_TLF_FIFO_blk[9] | proc_27_input_sync_blk[9] | proc_27_output_sync_blk[9]);
    assign proc_27_data_FIFO_blk[10] = 1'b0;
    assign proc_27_data_PIPO_blk[10] = 1'b0;
    assign proc_27_start_FIFO_blk[10] = 1'b0;
    assign proc_27_TLF_FIFO_blk[10] = 1'b0;
    assign proc_27_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_27_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_27[10] = dl_detect_out ? proc_dep_vld_vec_27_reg[10] : (proc_27_data_FIFO_blk[10] | proc_27_data_PIPO_blk[10] | proc_27_start_FIFO_blk[10] | proc_27_TLF_FIFO_blk[10] | proc_27_input_sync_blk[10] | proc_27_output_sync_blk[10]);
    assign proc_27_data_FIFO_blk[11] = 1'b0;
    assign proc_27_data_PIPO_blk[11] = 1'b0;
    assign proc_27_start_FIFO_blk[11] = 1'b0;
    assign proc_27_TLF_FIFO_blk[11] = 1'b0;
    assign proc_27_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_27_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_27[11] = dl_detect_out ? proc_dep_vld_vec_27_reg[11] : (proc_27_data_FIFO_blk[11] | proc_27_data_PIPO_blk[11] | proc_27_start_FIFO_blk[11] | proc_27_TLF_FIFO_blk[11] | proc_27_input_sync_blk[11] | proc_27_output_sync_blk[11]);
    assign proc_27_data_FIFO_blk[12] = 1'b0;
    assign proc_27_data_PIPO_blk[12] = 1'b0;
    assign proc_27_start_FIFO_blk[12] = 1'b0;
    assign proc_27_TLF_FIFO_blk[12] = 1'b0;
    assign proc_27_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_27_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_27[12] = dl_detect_out ? proc_dep_vld_vec_27_reg[12] : (proc_27_data_FIFO_blk[12] | proc_27_data_PIPO_blk[12] | proc_27_start_FIFO_blk[12] | proc_27_TLF_FIFO_blk[12] | proc_27_input_sync_blk[12] | proc_27_output_sync_blk[12]);
    assign proc_27_data_FIFO_blk[13] = 1'b0;
    assign proc_27_data_PIPO_blk[13] = 1'b0;
    assign proc_27_start_FIFO_blk[13] = 1'b0;
    assign proc_27_TLF_FIFO_blk[13] = 1'b0;
    assign proc_27_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_27_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_27[13] = dl_detect_out ? proc_dep_vld_vec_27_reg[13] : (proc_27_data_FIFO_blk[13] | proc_27_data_PIPO_blk[13] | proc_27_start_FIFO_blk[13] | proc_27_TLF_FIFO_blk[13] | proc_27_input_sync_blk[13] | proc_27_output_sync_blk[13]);
    assign proc_27_data_FIFO_blk[14] = 1'b0;
    assign proc_27_data_PIPO_blk[14] = 1'b0;
    assign proc_27_start_FIFO_blk[14] = 1'b0;
    assign proc_27_TLF_FIFO_blk[14] = 1'b0;
    assign proc_27_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_27_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_27[14] = dl_detect_out ? proc_dep_vld_vec_27_reg[14] : (proc_27_data_FIFO_blk[14] | proc_27_data_PIPO_blk[14] | proc_27_start_FIFO_blk[14] | proc_27_TLF_FIFO_blk[14] | proc_27_input_sync_blk[14] | proc_27_output_sync_blk[14]);
    assign proc_27_data_FIFO_blk[15] = 1'b0;
    assign proc_27_data_PIPO_blk[15] = 1'b0;
    assign proc_27_start_FIFO_blk[15] = 1'b0;
    assign proc_27_TLF_FIFO_blk[15] = 1'b0;
    assign proc_27_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_27_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_27[15] = dl_detect_out ? proc_dep_vld_vec_27_reg[15] : (proc_27_data_FIFO_blk[15] | proc_27_data_PIPO_blk[15] | proc_27_start_FIFO_blk[15] | proc_27_TLF_FIFO_blk[15] | proc_27_input_sync_blk[15] | proc_27_output_sync_blk[15]);
    assign proc_27_data_FIFO_blk[16] = 1'b0;
    assign proc_27_data_PIPO_blk[16] = 1'b0;
    assign proc_27_start_FIFO_blk[16] = 1'b0;
    assign proc_27_TLF_FIFO_blk[16] = 1'b0;
    assign proc_27_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_27_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_27[16] = dl_detect_out ? proc_dep_vld_vec_27_reg[16] : (proc_27_data_FIFO_blk[16] | proc_27_data_PIPO_blk[16] | proc_27_start_FIFO_blk[16] | proc_27_TLF_FIFO_blk[16] | proc_27_input_sync_blk[16] | proc_27_output_sync_blk[16]);
    assign proc_27_data_FIFO_blk[17] = 1'b0;
    assign proc_27_data_PIPO_blk[17] = 1'b0;
    assign proc_27_start_FIFO_blk[17] = 1'b0;
    assign proc_27_TLF_FIFO_blk[17] = 1'b0;
    assign proc_27_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_27_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_27[17] = dl_detect_out ? proc_dep_vld_vec_27_reg[17] : (proc_27_data_FIFO_blk[17] | proc_27_data_PIPO_blk[17] | proc_27_start_FIFO_blk[17] | proc_27_TLF_FIFO_blk[17] | proc_27_input_sync_blk[17] | proc_27_output_sync_blk[17]);
    assign proc_27_data_FIFO_blk[18] = 1'b0;
    assign proc_27_data_PIPO_blk[18] = 1'b0;
    assign proc_27_start_FIFO_blk[18] = 1'b0;
    assign proc_27_TLF_FIFO_blk[18] = 1'b0;
    assign proc_27_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_27_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_27[18] = dl_detect_out ? proc_dep_vld_vec_27_reg[18] : (proc_27_data_FIFO_blk[18] | proc_27_data_PIPO_blk[18] | proc_27_start_FIFO_blk[18] | proc_27_TLF_FIFO_blk[18] | proc_27_input_sync_blk[18] | proc_27_output_sync_blk[18]);
    assign proc_27_data_FIFO_blk[19] = 1'b0;
    assign proc_27_data_PIPO_blk[19] = 1'b0;
    assign proc_27_start_FIFO_blk[19] = 1'b0;
    assign proc_27_TLF_FIFO_blk[19] = 1'b0;
    assign proc_27_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_27_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_27[19] = dl_detect_out ? proc_dep_vld_vec_27_reg[19] : (proc_27_data_FIFO_blk[19] | proc_27_data_PIPO_blk[19] | proc_27_start_FIFO_blk[19] | proc_27_TLF_FIFO_blk[19] | proc_27_input_sync_blk[19] | proc_27_output_sync_blk[19]);
    assign proc_27_data_FIFO_blk[20] = 1'b0;
    assign proc_27_data_PIPO_blk[20] = 1'b0;
    assign proc_27_start_FIFO_blk[20] = 1'b0;
    assign proc_27_TLF_FIFO_blk[20] = 1'b0;
    assign proc_27_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_27_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_27[20] = dl_detect_out ? proc_dep_vld_vec_27_reg[20] : (proc_27_data_FIFO_blk[20] | proc_27_data_PIPO_blk[20] | proc_27_start_FIFO_blk[20] | proc_27_TLF_FIFO_blk[20] | proc_27_input_sync_blk[20] | proc_27_output_sync_blk[20]);
    assign proc_27_data_FIFO_blk[21] = 1'b0;
    assign proc_27_data_PIPO_blk[21] = 1'b0;
    assign proc_27_start_FIFO_blk[21] = 1'b0;
    assign proc_27_TLF_FIFO_blk[21] = 1'b0;
    assign proc_27_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_27_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_27[21] = dl_detect_out ? proc_dep_vld_vec_27_reg[21] : (proc_27_data_FIFO_blk[21] | proc_27_data_PIPO_blk[21] | proc_27_start_FIFO_blk[21] | proc_27_TLF_FIFO_blk[21] | proc_27_input_sync_blk[21] | proc_27_output_sync_blk[21]);
    assign proc_27_data_FIFO_blk[22] = 1'b0;
    assign proc_27_data_PIPO_blk[22] = 1'b0;
    assign proc_27_start_FIFO_blk[22] = 1'b0;
    assign proc_27_TLF_FIFO_blk[22] = 1'b0;
    assign proc_27_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_27_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_27[22] = dl_detect_out ? proc_dep_vld_vec_27_reg[22] : (proc_27_data_FIFO_blk[22] | proc_27_data_PIPO_blk[22] | proc_27_start_FIFO_blk[22] | proc_27_TLF_FIFO_blk[22] | proc_27_input_sync_blk[22] | proc_27_output_sync_blk[22]);
    assign proc_27_data_FIFO_blk[23] = 1'b0;
    assign proc_27_data_PIPO_blk[23] = 1'b0;
    assign proc_27_start_FIFO_blk[23] = 1'b0;
    assign proc_27_TLF_FIFO_blk[23] = 1'b0;
    assign proc_27_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_27_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_27[23] = dl_detect_out ? proc_dep_vld_vec_27_reg[23] : (proc_27_data_FIFO_blk[23] | proc_27_data_PIPO_blk[23] | proc_27_start_FIFO_blk[23] | proc_27_TLF_FIFO_blk[23] | proc_27_input_sync_blk[23] | proc_27_output_sync_blk[23]);
    assign proc_27_data_FIFO_blk[24] = 1'b0;
    assign proc_27_data_PIPO_blk[24] = 1'b0;
    assign proc_27_start_FIFO_blk[24] = 1'b0;
    assign proc_27_TLF_FIFO_blk[24] = 1'b0;
    assign proc_27_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_27_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_27[24] = dl_detect_out ? proc_dep_vld_vec_27_reg[24] : (proc_27_data_FIFO_blk[24] | proc_27_data_PIPO_blk[24] | proc_27_start_FIFO_blk[24] | proc_27_TLF_FIFO_blk[24] | proc_27_input_sync_blk[24] | proc_27_output_sync_blk[24]);
    assign proc_27_data_FIFO_blk[25] = 1'b0;
    assign proc_27_data_PIPO_blk[25] = 1'b0;
    assign proc_27_start_FIFO_blk[25] = 1'b0;
    assign proc_27_TLF_FIFO_blk[25] = 1'b0;
    assign proc_27_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_27_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_27[25] = dl_detect_out ? proc_dep_vld_vec_27_reg[25] : (proc_27_data_FIFO_blk[25] | proc_27_data_PIPO_blk[25] | proc_27_start_FIFO_blk[25] | proc_27_TLF_FIFO_blk[25] | proc_27_input_sync_blk[25] | proc_27_output_sync_blk[25]);
    assign proc_27_data_FIFO_blk[26] = 1'b0;
    assign proc_27_data_PIPO_blk[26] = 1'b0;
    assign proc_27_start_FIFO_blk[26] = 1'b0;
    assign proc_27_TLF_FIFO_blk[26] = 1'b0;
    assign proc_27_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_27_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_27[26] = dl_detect_out ? proc_dep_vld_vec_27_reg[26] : (proc_27_data_FIFO_blk[26] | proc_27_data_PIPO_blk[26] | proc_27_start_FIFO_blk[26] | proc_27_TLF_FIFO_blk[26] | proc_27_input_sync_blk[26] | proc_27_output_sync_blk[26]);
    assign proc_27_data_FIFO_blk[27] = 1'b0;
    assign proc_27_data_PIPO_blk[27] = 1'b0;
    assign proc_27_start_FIFO_blk[27] = 1'b0;
    assign proc_27_TLF_FIFO_blk[27] = 1'b0;
    assign proc_27_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_27_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_27[27] = dl_detect_out ? proc_dep_vld_vec_27_reg[27] : (proc_27_data_FIFO_blk[27] | proc_27_data_PIPO_blk[27] | proc_27_start_FIFO_blk[27] | proc_27_TLF_FIFO_blk[27] | proc_27_input_sync_blk[27] | proc_27_output_sync_blk[27]);
    assign proc_27_data_FIFO_blk[28] = 1'b0;
    assign proc_27_data_PIPO_blk[28] = 1'b0;
    assign proc_27_start_FIFO_blk[28] = 1'b0;
    assign proc_27_TLF_FIFO_blk[28] = 1'b0;
    assign proc_27_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_27_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_27[28] = dl_detect_out ? proc_dep_vld_vec_27_reg[28] : (proc_27_data_FIFO_blk[28] | proc_27_data_PIPO_blk[28] | proc_27_start_FIFO_blk[28] | proc_27_TLF_FIFO_blk[28] | proc_27_input_sync_blk[28] | proc_27_output_sync_blk[28]);
    assign proc_27_data_FIFO_blk[29] = 1'b0;
    assign proc_27_data_PIPO_blk[29] = 1'b0;
    assign proc_27_start_FIFO_blk[29] = 1'b0;
    assign proc_27_TLF_FIFO_blk[29] = 1'b0;
    assign proc_27_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_27_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_27[29] = dl_detect_out ? proc_dep_vld_vec_27_reg[29] : (proc_27_data_FIFO_blk[29] | proc_27_data_PIPO_blk[29] | proc_27_start_FIFO_blk[29] | proc_27_TLF_FIFO_blk[29] | proc_27_input_sync_blk[29] | proc_27_output_sync_blk[29]);
    assign proc_27_data_FIFO_blk[30] = 1'b0;
    assign proc_27_data_PIPO_blk[30] = 1'b0;
    assign proc_27_start_FIFO_blk[30] = 1'b0;
    assign proc_27_TLF_FIFO_blk[30] = 1'b0;
    assign proc_27_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_27_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_27[30] = dl_detect_out ? proc_dep_vld_vec_27_reg[30] : (proc_27_data_FIFO_blk[30] | proc_27_data_PIPO_blk[30] | proc_27_start_FIFO_blk[30] | proc_27_TLF_FIFO_blk[30] | proc_27_input_sync_blk[30] | proc_27_output_sync_blk[30]);
    assign proc_27_data_FIFO_blk[31] = 1'b0;
    assign proc_27_data_PIPO_blk[31] = 1'b0;
    assign proc_27_start_FIFO_blk[31] = 1'b0;
    assign proc_27_TLF_FIFO_blk[31] = 1'b0;
    assign proc_27_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_27_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_27[31] = dl_detect_out ? proc_dep_vld_vec_27_reg[31] : (proc_27_data_FIFO_blk[31] | proc_27_data_PIPO_blk[31] | proc_27_start_FIFO_blk[31] | proc_27_TLF_FIFO_blk[31] | proc_27_input_sync_blk[31] | proc_27_output_sync_blk[31]);
    assign proc_27_data_FIFO_blk[32] = 1'b0;
    assign proc_27_data_PIPO_blk[32] = 1'b0;
    assign proc_27_start_FIFO_blk[32] = 1'b0;
    assign proc_27_TLF_FIFO_blk[32] = 1'b0;
    assign proc_27_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_22_U0_ap_ready & ProcessingElement_22_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_27_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_27[32] = dl_detect_out ? proc_dep_vld_vec_27_reg[32] : (proc_27_data_FIFO_blk[32] | proc_27_data_PIPO_blk[32] | proc_27_start_FIFO_blk[32] | proc_27_TLF_FIFO_blk[32] | proc_27_input_sync_blk[32] | proc_27_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_27_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_27_reg <= proc_dep_vld_vec_27;
        end
    end
    assign in_chan_dep_vld_vec_27[0] = dep_chan_vld_0_27;
    assign in_chan_dep_data_vec_27[39 : 0] = dep_chan_data_0_27;
    assign token_in_vec_27[0] = token_0_27;
    assign in_chan_dep_vld_vec_27[1] = dep_chan_vld_1_27;
    assign in_chan_dep_data_vec_27[79 : 40] = dep_chan_data_1_27;
    assign token_in_vec_27[1] = token_1_27;
    assign in_chan_dep_vld_vec_27[2] = dep_chan_vld_3_27;
    assign in_chan_dep_data_vec_27[119 : 80] = dep_chan_data_3_27;
    assign token_in_vec_27[2] = token_3_27;
    assign in_chan_dep_vld_vec_27[3] = dep_chan_vld_6_27;
    assign in_chan_dep_data_vec_27[159 : 120] = dep_chan_data_6_27;
    assign token_in_vec_27[3] = token_6_27;
    assign in_chan_dep_vld_vec_27[4] = dep_chan_vld_7_27;
    assign in_chan_dep_data_vec_27[199 : 160] = dep_chan_data_7_27;
    assign token_in_vec_27[4] = token_7_27;
    assign in_chan_dep_vld_vec_27[5] = dep_chan_vld_8_27;
    assign in_chan_dep_data_vec_27[239 : 200] = dep_chan_data_8_27;
    assign token_in_vec_27[5] = token_8_27;
    assign in_chan_dep_vld_vec_27[6] = dep_chan_vld_9_27;
    assign in_chan_dep_data_vec_27[279 : 240] = dep_chan_data_9_27;
    assign token_in_vec_27[6] = token_9_27;
    assign in_chan_dep_vld_vec_27[7] = dep_chan_vld_10_27;
    assign in_chan_dep_data_vec_27[319 : 280] = dep_chan_data_10_27;
    assign token_in_vec_27[7] = token_10_27;
    assign in_chan_dep_vld_vec_27[8] = dep_chan_vld_11_27;
    assign in_chan_dep_data_vec_27[359 : 320] = dep_chan_data_11_27;
    assign token_in_vec_27[8] = token_11_27;
    assign in_chan_dep_vld_vec_27[9] = dep_chan_vld_12_27;
    assign in_chan_dep_data_vec_27[399 : 360] = dep_chan_data_12_27;
    assign token_in_vec_27[9] = token_12_27;
    assign in_chan_dep_vld_vec_27[10] = dep_chan_vld_13_27;
    assign in_chan_dep_data_vec_27[439 : 400] = dep_chan_data_13_27;
    assign token_in_vec_27[10] = token_13_27;
    assign in_chan_dep_vld_vec_27[11] = dep_chan_vld_14_27;
    assign in_chan_dep_data_vec_27[479 : 440] = dep_chan_data_14_27;
    assign token_in_vec_27[11] = token_14_27;
    assign in_chan_dep_vld_vec_27[12] = dep_chan_vld_15_27;
    assign in_chan_dep_data_vec_27[519 : 480] = dep_chan_data_15_27;
    assign token_in_vec_27[12] = token_15_27;
    assign in_chan_dep_vld_vec_27[13] = dep_chan_vld_16_27;
    assign in_chan_dep_data_vec_27[559 : 520] = dep_chan_data_16_27;
    assign token_in_vec_27[13] = token_16_27;
    assign in_chan_dep_vld_vec_27[14] = dep_chan_vld_17_27;
    assign in_chan_dep_data_vec_27[599 : 560] = dep_chan_data_17_27;
    assign token_in_vec_27[14] = token_17_27;
    assign in_chan_dep_vld_vec_27[15] = dep_chan_vld_18_27;
    assign in_chan_dep_data_vec_27[639 : 600] = dep_chan_data_18_27;
    assign token_in_vec_27[15] = token_18_27;
    assign in_chan_dep_vld_vec_27[16] = dep_chan_vld_19_27;
    assign in_chan_dep_data_vec_27[679 : 640] = dep_chan_data_19_27;
    assign token_in_vec_27[16] = token_19_27;
    assign in_chan_dep_vld_vec_27[17] = dep_chan_vld_20_27;
    assign in_chan_dep_data_vec_27[719 : 680] = dep_chan_data_20_27;
    assign token_in_vec_27[17] = token_20_27;
    assign in_chan_dep_vld_vec_27[18] = dep_chan_vld_21_27;
    assign in_chan_dep_data_vec_27[759 : 720] = dep_chan_data_21_27;
    assign token_in_vec_27[18] = token_21_27;
    assign in_chan_dep_vld_vec_27[19] = dep_chan_vld_22_27;
    assign in_chan_dep_data_vec_27[799 : 760] = dep_chan_data_22_27;
    assign token_in_vec_27[19] = token_22_27;
    assign in_chan_dep_vld_vec_27[20] = dep_chan_vld_23_27;
    assign in_chan_dep_data_vec_27[839 : 800] = dep_chan_data_23_27;
    assign token_in_vec_27[20] = token_23_27;
    assign in_chan_dep_vld_vec_27[21] = dep_chan_vld_24_27;
    assign in_chan_dep_data_vec_27[879 : 840] = dep_chan_data_24_27;
    assign token_in_vec_27[21] = token_24_27;
    assign in_chan_dep_vld_vec_27[22] = dep_chan_vld_25_27;
    assign in_chan_dep_data_vec_27[919 : 880] = dep_chan_data_25_27;
    assign token_in_vec_27[22] = token_25_27;
    assign in_chan_dep_vld_vec_27[23] = dep_chan_vld_26_27;
    assign in_chan_dep_data_vec_27[959 : 920] = dep_chan_data_26_27;
    assign token_in_vec_27[23] = token_26_27;
    assign in_chan_dep_vld_vec_27[24] = dep_chan_vld_28_27;
    assign in_chan_dep_data_vec_27[999 : 960] = dep_chan_data_28_27;
    assign token_in_vec_27[24] = token_28_27;
    assign in_chan_dep_vld_vec_27[25] = dep_chan_vld_29_27;
    assign in_chan_dep_data_vec_27[1039 : 1000] = dep_chan_data_29_27;
    assign token_in_vec_27[25] = token_29_27;
    assign in_chan_dep_vld_vec_27[26] = dep_chan_vld_30_27;
    assign in_chan_dep_data_vec_27[1079 : 1040] = dep_chan_data_30_27;
    assign token_in_vec_27[26] = token_30_27;
    assign in_chan_dep_vld_vec_27[27] = dep_chan_vld_31_27;
    assign in_chan_dep_data_vec_27[1119 : 1080] = dep_chan_data_31_27;
    assign token_in_vec_27[27] = token_31_27;
    assign in_chan_dep_vld_vec_27[28] = dep_chan_vld_32_27;
    assign in_chan_dep_data_vec_27[1159 : 1120] = dep_chan_data_32_27;
    assign token_in_vec_27[28] = token_32_27;
    assign in_chan_dep_vld_vec_27[29] = dep_chan_vld_33_27;
    assign in_chan_dep_data_vec_27[1199 : 1160] = dep_chan_data_33_27;
    assign token_in_vec_27[29] = token_33_27;
    assign in_chan_dep_vld_vec_27[30] = dep_chan_vld_34_27;
    assign in_chan_dep_data_vec_27[1239 : 1200] = dep_chan_data_34_27;
    assign token_in_vec_27[30] = token_34_27;
    assign in_chan_dep_vld_vec_27[31] = dep_chan_vld_35_27;
    assign in_chan_dep_data_vec_27[1279 : 1240] = dep_chan_data_35_27;
    assign token_in_vec_27[31] = token_35_27;
    assign in_chan_dep_vld_vec_27[32] = dep_chan_vld_36_27;
    assign in_chan_dep_data_vec_27[1319 : 1280] = dep_chan_data_36_27;
    assign token_in_vec_27[32] = token_36_27;
    assign dep_chan_vld_27_26 = out_chan_dep_vld_vec_27[0];
    assign dep_chan_data_27_26 = out_chan_dep_data_27;
    assign token_27_26 = token_out_vec_27[0];
    assign dep_chan_vld_27_28 = out_chan_dep_vld_vec_27[1];
    assign dep_chan_data_27_28 = out_chan_dep_data_27;
    assign token_27_28 = token_out_vec_27[1];
    assign dep_chan_vld_27_0 = out_chan_dep_vld_vec_27[2];
    assign dep_chan_data_27_0 = out_chan_dep_data_27;
    assign token_27_0 = token_out_vec_27[2];
    assign dep_chan_vld_27_1 = out_chan_dep_vld_vec_27[3];
    assign dep_chan_data_27_1 = out_chan_dep_data_27;
    assign token_27_1 = token_out_vec_27[3];
    assign dep_chan_vld_27_3 = out_chan_dep_vld_vec_27[4];
    assign dep_chan_data_27_3 = out_chan_dep_data_27;
    assign token_27_3 = token_out_vec_27[4];
    assign dep_chan_vld_27_6 = out_chan_dep_vld_vec_27[5];
    assign dep_chan_data_27_6 = out_chan_dep_data_27;
    assign token_27_6 = token_out_vec_27[5];
    assign dep_chan_vld_27_7 = out_chan_dep_vld_vec_27[6];
    assign dep_chan_data_27_7 = out_chan_dep_data_27;
    assign token_27_7 = token_out_vec_27[6];
    assign dep_chan_vld_27_8 = out_chan_dep_vld_vec_27[7];
    assign dep_chan_data_27_8 = out_chan_dep_data_27;
    assign token_27_8 = token_out_vec_27[7];
    assign dep_chan_vld_27_9 = out_chan_dep_vld_vec_27[8];
    assign dep_chan_data_27_9 = out_chan_dep_data_27;
    assign token_27_9 = token_out_vec_27[8];
    assign dep_chan_vld_27_10 = out_chan_dep_vld_vec_27[9];
    assign dep_chan_data_27_10 = out_chan_dep_data_27;
    assign token_27_10 = token_out_vec_27[9];
    assign dep_chan_vld_27_11 = out_chan_dep_vld_vec_27[10];
    assign dep_chan_data_27_11 = out_chan_dep_data_27;
    assign token_27_11 = token_out_vec_27[10];
    assign dep_chan_vld_27_12 = out_chan_dep_vld_vec_27[11];
    assign dep_chan_data_27_12 = out_chan_dep_data_27;
    assign token_27_12 = token_out_vec_27[11];
    assign dep_chan_vld_27_13 = out_chan_dep_vld_vec_27[12];
    assign dep_chan_data_27_13 = out_chan_dep_data_27;
    assign token_27_13 = token_out_vec_27[12];
    assign dep_chan_vld_27_14 = out_chan_dep_vld_vec_27[13];
    assign dep_chan_data_27_14 = out_chan_dep_data_27;
    assign token_27_14 = token_out_vec_27[13];
    assign dep_chan_vld_27_15 = out_chan_dep_vld_vec_27[14];
    assign dep_chan_data_27_15 = out_chan_dep_data_27;
    assign token_27_15 = token_out_vec_27[14];
    assign dep_chan_vld_27_16 = out_chan_dep_vld_vec_27[15];
    assign dep_chan_data_27_16 = out_chan_dep_data_27;
    assign token_27_16 = token_out_vec_27[15];
    assign dep_chan_vld_27_17 = out_chan_dep_vld_vec_27[16];
    assign dep_chan_data_27_17 = out_chan_dep_data_27;
    assign token_27_17 = token_out_vec_27[16];
    assign dep_chan_vld_27_18 = out_chan_dep_vld_vec_27[17];
    assign dep_chan_data_27_18 = out_chan_dep_data_27;
    assign token_27_18 = token_out_vec_27[17];
    assign dep_chan_vld_27_19 = out_chan_dep_vld_vec_27[18];
    assign dep_chan_data_27_19 = out_chan_dep_data_27;
    assign token_27_19 = token_out_vec_27[18];
    assign dep_chan_vld_27_20 = out_chan_dep_vld_vec_27[19];
    assign dep_chan_data_27_20 = out_chan_dep_data_27;
    assign token_27_20 = token_out_vec_27[19];
    assign dep_chan_vld_27_21 = out_chan_dep_vld_vec_27[20];
    assign dep_chan_data_27_21 = out_chan_dep_data_27;
    assign token_27_21 = token_out_vec_27[20];
    assign dep_chan_vld_27_22 = out_chan_dep_vld_vec_27[21];
    assign dep_chan_data_27_22 = out_chan_dep_data_27;
    assign token_27_22 = token_out_vec_27[21];
    assign dep_chan_vld_27_23 = out_chan_dep_vld_vec_27[22];
    assign dep_chan_data_27_23 = out_chan_dep_data_27;
    assign token_27_23 = token_out_vec_27[22];
    assign dep_chan_vld_27_24 = out_chan_dep_vld_vec_27[23];
    assign dep_chan_data_27_24 = out_chan_dep_data_27;
    assign token_27_24 = token_out_vec_27[23];
    assign dep_chan_vld_27_25 = out_chan_dep_vld_vec_27[24];
    assign dep_chan_data_27_25 = out_chan_dep_data_27;
    assign token_27_25 = token_out_vec_27[24];
    assign dep_chan_vld_27_29 = out_chan_dep_vld_vec_27[25];
    assign dep_chan_data_27_29 = out_chan_dep_data_27;
    assign token_27_29 = token_out_vec_27[25];
    assign dep_chan_vld_27_30 = out_chan_dep_vld_vec_27[26];
    assign dep_chan_data_27_30 = out_chan_dep_data_27;
    assign token_27_30 = token_out_vec_27[26];
    assign dep_chan_vld_27_31 = out_chan_dep_vld_vec_27[27];
    assign dep_chan_data_27_31 = out_chan_dep_data_27;
    assign token_27_31 = token_out_vec_27[27];
    assign dep_chan_vld_27_32 = out_chan_dep_vld_vec_27[28];
    assign dep_chan_data_27_32 = out_chan_dep_data_27;
    assign token_27_32 = token_out_vec_27[28];
    assign dep_chan_vld_27_33 = out_chan_dep_vld_vec_27[29];
    assign dep_chan_data_27_33 = out_chan_dep_data_27;
    assign token_27_33 = token_out_vec_27[29];
    assign dep_chan_vld_27_34 = out_chan_dep_vld_vec_27[30];
    assign dep_chan_data_27_34 = out_chan_dep_data_27;
    assign token_27_34 = token_out_vec_27[30];
    assign dep_chan_vld_27_35 = out_chan_dep_vld_vec_27[31];
    assign dep_chan_data_27_35 = out_chan_dep_data_27;
    assign token_27_35 = token_out_vec_27[31];
    assign dep_chan_vld_27_36 = out_chan_dep_vld_vec_27[32];
    assign dep_chan_data_27_36 = out_chan_dep_data_27;
    assign token_27_36 = token_out_vec_27[32];

    // Process: ProcessingElement_23_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 28, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_28 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_28),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_28),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_28),
        .token_in_vec(token_in_vec_28),
        .dl_detect_in(dl_detect_out),
        .origin(origin[28]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_28),
        .out_chan_dep_data(out_chan_dep_data_28),
        .token_out_vec(token_out_vec_28),
        .dl_detect_out(dl_in_vec[28]));

    assign proc_28_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_22_blk_n) | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_22_blk_n) | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_WriteC_Flattened_fu_179.cPipes_22_blk_n);
    assign proc_28_data_PIPO_blk[0] = 1'b0;
    assign proc_28_start_FIFO_blk[0] = 1'b0;
    assign proc_28_TLF_FIFO_blk[0] = 1'b0;
    assign proc_28_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_28_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_28[0] = dl_detect_out ? proc_dep_vld_vec_28_reg[0] : (proc_28_data_FIFO_blk[0] | proc_28_data_PIPO_blk[0] | proc_28_start_FIFO_blk[0] | proc_28_TLF_FIFO_blk[0] | proc_28_input_sync_blk[0] | proc_28_output_sync_blk[0]);
    assign proc_28_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_23_blk_n) | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_23_blk_n) | (~ProcessingElement_23_U0.grp_ProcessingElement_23_Pipeline_WriteC_Flattened_fu_179.cPipes_23_blk_n);
    assign proc_28_data_PIPO_blk[1] = 1'b0;
    assign proc_28_start_FIFO_blk[1] = 1'b0;
    assign proc_28_TLF_FIFO_blk[1] = 1'b0;
    assign proc_28_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_28_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_28[1] = dl_detect_out ? proc_dep_vld_vec_28_reg[1] : (proc_28_data_FIFO_blk[1] | proc_28_data_PIPO_blk[1] | proc_28_start_FIFO_blk[1] | proc_28_TLF_FIFO_blk[1] | proc_28_input_sync_blk[1] | proc_28_output_sync_blk[1]);
    assign proc_28_data_FIFO_blk[2] = 1'b0;
    assign proc_28_data_PIPO_blk[2] = 1'b0;
    assign proc_28_start_FIFO_blk[2] = 1'b0;
    assign proc_28_TLF_FIFO_blk[2] = 1'b0;
    assign proc_28_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_28_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_28[2] = dl_detect_out ? proc_dep_vld_vec_28_reg[2] : (proc_28_data_FIFO_blk[2] | proc_28_data_PIPO_blk[2] | proc_28_start_FIFO_blk[2] | proc_28_TLF_FIFO_blk[2] | proc_28_input_sync_blk[2] | proc_28_output_sync_blk[2]);
    assign proc_28_data_FIFO_blk[3] = 1'b0;
    assign proc_28_data_PIPO_blk[3] = 1'b0;
    assign proc_28_start_FIFO_blk[3] = 1'b0;
    assign proc_28_TLF_FIFO_blk[3] = 1'b0;
    assign proc_28_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_28_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_28[3] = dl_detect_out ? proc_dep_vld_vec_28_reg[3] : (proc_28_data_FIFO_blk[3] | proc_28_data_PIPO_blk[3] | proc_28_start_FIFO_blk[3] | proc_28_TLF_FIFO_blk[3] | proc_28_input_sync_blk[3] | proc_28_output_sync_blk[3]);
    assign proc_28_data_FIFO_blk[4] = 1'b0;
    assign proc_28_data_PIPO_blk[4] = 1'b0;
    assign proc_28_start_FIFO_blk[4] = 1'b0;
    assign proc_28_TLF_FIFO_blk[4] = 1'b0;
    assign proc_28_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_28_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_28[4] = dl_detect_out ? proc_dep_vld_vec_28_reg[4] : (proc_28_data_FIFO_blk[4] | proc_28_data_PIPO_blk[4] | proc_28_start_FIFO_blk[4] | proc_28_TLF_FIFO_blk[4] | proc_28_input_sync_blk[4] | proc_28_output_sync_blk[4]);
    assign proc_28_data_FIFO_blk[5] = 1'b0;
    assign proc_28_data_PIPO_blk[5] = 1'b0;
    assign proc_28_start_FIFO_blk[5] = 1'b0;
    assign proc_28_TLF_FIFO_blk[5] = 1'b0;
    assign proc_28_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_28_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_28[5] = dl_detect_out ? proc_dep_vld_vec_28_reg[5] : (proc_28_data_FIFO_blk[5] | proc_28_data_PIPO_blk[5] | proc_28_start_FIFO_blk[5] | proc_28_TLF_FIFO_blk[5] | proc_28_input_sync_blk[5] | proc_28_output_sync_blk[5]);
    assign proc_28_data_FIFO_blk[6] = 1'b0;
    assign proc_28_data_PIPO_blk[6] = 1'b0;
    assign proc_28_start_FIFO_blk[6] = 1'b0;
    assign proc_28_TLF_FIFO_blk[6] = 1'b0;
    assign proc_28_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_28_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_28[6] = dl_detect_out ? proc_dep_vld_vec_28_reg[6] : (proc_28_data_FIFO_blk[6] | proc_28_data_PIPO_blk[6] | proc_28_start_FIFO_blk[6] | proc_28_TLF_FIFO_blk[6] | proc_28_input_sync_blk[6] | proc_28_output_sync_blk[6]);
    assign proc_28_data_FIFO_blk[7] = 1'b0;
    assign proc_28_data_PIPO_blk[7] = 1'b0;
    assign proc_28_start_FIFO_blk[7] = 1'b0;
    assign proc_28_TLF_FIFO_blk[7] = 1'b0;
    assign proc_28_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_28_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_28[7] = dl_detect_out ? proc_dep_vld_vec_28_reg[7] : (proc_28_data_FIFO_blk[7] | proc_28_data_PIPO_blk[7] | proc_28_start_FIFO_blk[7] | proc_28_TLF_FIFO_blk[7] | proc_28_input_sync_blk[7] | proc_28_output_sync_blk[7]);
    assign proc_28_data_FIFO_blk[8] = 1'b0;
    assign proc_28_data_PIPO_blk[8] = 1'b0;
    assign proc_28_start_FIFO_blk[8] = 1'b0;
    assign proc_28_TLF_FIFO_blk[8] = 1'b0;
    assign proc_28_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_28_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_28[8] = dl_detect_out ? proc_dep_vld_vec_28_reg[8] : (proc_28_data_FIFO_blk[8] | proc_28_data_PIPO_blk[8] | proc_28_start_FIFO_blk[8] | proc_28_TLF_FIFO_blk[8] | proc_28_input_sync_blk[8] | proc_28_output_sync_blk[8]);
    assign proc_28_data_FIFO_blk[9] = 1'b0;
    assign proc_28_data_PIPO_blk[9] = 1'b0;
    assign proc_28_start_FIFO_blk[9] = 1'b0;
    assign proc_28_TLF_FIFO_blk[9] = 1'b0;
    assign proc_28_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_28_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_28[9] = dl_detect_out ? proc_dep_vld_vec_28_reg[9] : (proc_28_data_FIFO_blk[9] | proc_28_data_PIPO_blk[9] | proc_28_start_FIFO_blk[9] | proc_28_TLF_FIFO_blk[9] | proc_28_input_sync_blk[9] | proc_28_output_sync_blk[9]);
    assign proc_28_data_FIFO_blk[10] = 1'b0;
    assign proc_28_data_PIPO_blk[10] = 1'b0;
    assign proc_28_start_FIFO_blk[10] = 1'b0;
    assign proc_28_TLF_FIFO_blk[10] = 1'b0;
    assign proc_28_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_28_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_28[10] = dl_detect_out ? proc_dep_vld_vec_28_reg[10] : (proc_28_data_FIFO_blk[10] | proc_28_data_PIPO_blk[10] | proc_28_start_FIFO_blk[10] | proc_28_TLF_FIFO_blk[10] | proc_28_input_sync_blk[10] | proc_28_output_sync_blk[10]);
    assign proc_28_data_FIFO_blk[11] = 1'b0;
    assign proc_28_data_PIPO_blk[11] = 1'b0;
    assign proc_28_start_FIFO_blk[11] = 1'b0;
    assign proc_28_TLF_FIFO_blk[11] = 1'b0;
    assign proc_28_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_28_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_28[11] = dl_detect_out ? proc_dep_vld_vec_28_reg[11] : (proc_28_data_FIFO_blk[11] | proc_28_data_PIPO_blk[11] | proc_28_start_FIFO_blk[11] | proc_28_TLF_FIFO_blk[11] | proc_28_input_sync_blk[11] | proc_28_output_sync_blk[11]);
    assign proc_28_data_FIFO_blk[12] = 1'b0;
    assign proc_28_data_PIPO_blk[12] = 1'b0;
    assign proc_28_start_FIFO_blk[12] = 1'b0;
    assign proc_28_TLF_FIFO_blk[12] = 1'b0;
    assign proc_28_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_28_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_28[12] = dl_detect_out ? proc_dep_vld_vec_28_reg[12] : (proc_28_data_FIFO_blk[12] | proc_28_data_PIPO_blk[12] | proc_28_start_FIFO_blk[12] | proc_28_TLF_FIFO_blk[12] | proc_28_input_sync_blk[12] | proc_28_output_sync_blk[12]);
    assign proc_28_data_FIFO_blk[13] = 1'b0;
    assign proc_28_data_PIPO_blk[13] = 1'b0;
    assign proc_28_start_FIFO_blk[13] = 1'b0;
    assign proc_28_TLF_FIFO_blk[13] = 1'b0;
    assign proc_28_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_28_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_28[13] = dl_detect_out ? proc_dep_vld_vec_28_reg[13] : (proc_28_data_FIFO_blk[13] | proc_28_data_PIPO_blk[13] | proc_28_start_FIFO_blk[13] | proc_28_TLF_FIFO_blk[13] | proc_28_input_sync_blk[13] | proc_28_output_sync_blk[13]);
    assign proc_28_data_FIFO_blk[14] = 1'b0;
    assign proc_28_data_PIPO_blk[14] = 1'b0;
    assign proc_28_start_FIFO_blk[14] = 1'b0;
    assign proc_28_TLF_FIFO_blk[14] = 1'b0;
    assign proc_28_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_28_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_28[14] = dl_detect_out ? proc_dep_vld_vec_28_reg[14] : (proc_28_data_FIFO_blk[14] | proc_28_data_PIPO_blk[14] | proc_28_start_FIFO_blk[14] | proc_28_TLF_FIFO_blk[14] | proc_28_input_sync_blk[14] | proc_28_output_sync_blk[14]);
    assign proc_28_data_FIFO_blk[15] = 1'b0;
    assign proc_28_data_PIPO_blk[15] = 1'b0;
    assign proc_28_start_FIFO_blk[15] = 1'b0;
    assign proc_28_TLF_FIFO_blk[15] = 1'b0;
    assign proc_28_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_28_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_28[15] = dl_detect_out ? proc_dep_vld_vec_28_reg[15] : (proc_28_data_FIFO_blk[15] | proc_28_data_PIPO_blk[15] | proc_28_start_FIFO_blk[15] | proc_28_TLF_FIFO_blk[15] | proc_28_input_sync_blk[15] | proc_28_output_sync_blk[15]);
    assign proc_28_data_FIFO_blk[16] = 1'b0;
    assign proc_28_data_PIPO_blk[16] = 1'b0;
    assign proc_28_start_FIFO_blk[16] = 1'b0;
    assign proc_28_TLF_FIFO_blk[16] = 1'b0;
    assign proc_28_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_28_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_28[16] = dl_detect_out ? proc_dep_vld_vec_28_reg[16] : (proc_28_data_FIFO_blk[16] | proc_28_data_PIPO_blk[16] | proc_28_start_FIFO_blk[16] | proc_28_TLF_FIFO_blk[16] | proc_28_input_sync_blk[16] | proc_28_output_sync_blk[16]);
    assign proc_28_data_FIFO_blk[17] = 1'b0;
    assign proc_28_data_PIPO_blk[17] = 1'b0;
    assign proc_28_start_FIFO_blk[17] = 1'b0;
    assign proc_28_TLF_FIFO_blk[17] = 1'b0;
    assign proc_28_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_28_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_28[17] = dl_detect_out ? proc_dep_vld_vec_28_reg[17] : (proc_28_data_FIFO_blk[17] | proc_28_data_PIPO_blk[17] | proc_28_start_FIFO_blk[17] | proc_28_TLF_FIFO_blk[17] | proc_28_input_sync_blk[17] | proc_28_output_sync_blk[17]);
    assign proc_28_data_FIFO_blk[18] = 1'b0;
    assign proc_28_data_PIPO_blk[18] = 1'b0;
    assign proc_28_start_FIFO_blk[18] = 1'b0;
    assign proc_28_TLF_FIFO_blk[18] = 1'b0;
    assign proc_28_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_28_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_28[18] = dl_detect_out ? proc_dep_vld_vec_28_reg[18] : (proc_28_data_FIFO_blk[18] | proc_28_data_PIPO_blk[18] | proc_28_start_FIFO_blk[18] | proc_28_TLF_FIFO_blk[18] | proc_28_input_sync_blk[18] | proc_28_output_sync_blk[18]);
    assign proc_28_data_FIFO_blk[19] = 1'b0;
    assign proc_28_data_PIPO_blk[19] = 1'b0;
    assign proc_28_start_FIFO_blk[19] = 1'b0;
    assign proc_28_TLF_FIFO_blk[19] = 1'b0;
    assign proc_28_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_28_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_28[19] = dl_detect_out ? proc_dep_vld_vec_28_reg[19] : (proc_28_data_FIFO_blk[19] | proc_28_data_PIPO_blk[19] | proc_28_start_FIFO_blk[19] | proc_28_TLF_FIFO_blk[19] | proc_28_input_sync_blk[19] | proc_28_output_sync_blk[19]);
    assign proc_28_data_FIFO_blk[20] = 1'b0;
    assign proc_28_data_PIPO_blk[20] = 1'b0;
    assign proc_28_start_FIFO_blk[20] = 1'b0;
    assign proc_28_TLF_FIFO_blk[20] = 1'b0;
    assign proc_28_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_28_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_28[20] = dl_detect_out ? proc_dep_vld_vec_28_reg[20] : (proc_28_data_FIFO_blk[20] | proc_28_data_PIPO_blk[20] | proc_28_start_FIFO_blk[20] | proc_28_TLF_FIFO_blk[20] | proc_28_input_sync_blk[20] | proc_28_output_sync_blk[20]);
    assign proc_28_data_FIFO_blk[21] = 1'b0;
    assign proc_28_data_PIPO_blk[21] = 1'b0;
    assign proc_28_start_FIFO_blk[21] = 1'b0;
    assign proc_28_TLF_FIFO_blk[21] = 1'b0;
    assign proc_28_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_28_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_28[21] = dl_detect_out ? proc_dep_vld_vec_28_reg[21] : (proc_28_data_FIFO_blk[21] | proc_28_data_PIPO_blk[21] | proc_28_start_FIFO_blk[21] | proc_28_TLF_FIFO_blk[21] | proc_28_input_sync_blk[21] | proc_28_output_sync_blk[21]);
    assign proc_28_data_FIFO_blk[22] = 1'b0;
    assign proc_28_data_PIPO_blk[22] = 1'b0;
    assign proc_28_start_FIFO_blk[22] = 1'b0;
    assign proc_28_TLF_FIFO_blk[22] = 1'b0;
    assign proc_28_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_28_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_28[22] = dl_detect_out ? proc_dep_vld_vec_28_reg[22] : (proc_28_data_FIFO_blk[22] | proc_28_data_PIPO_blk[22] | proc_28_start_FIFO_blk[22] | proc_28_TLF_FIFO_blk[22] | proc_28_input_sync_blk[22] | proc_28_output_sync_blk[22]);
    assign proc_28_data_FIFO_blk[23] = 1'b0;
    assign proc_28_data_PIPO_blk[23] = 1'b0;
    assign proc_28_start_FIFO_blk[23] = 1'b0;
    assign proc_28_TLF_FIFO_blk[23] = 1'b0;
    assign proc_28_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_28_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_28[23] = dl_detect_out ? proc_dep_vld_vec_28_reg[23] : (proc_28_data_FIFO_blk[23] | proc_28_data_PIPO_blk[23] | proc_28_start_FIFO_blk[23] | proc_28_TLF_FIFO_blk[23] | proc_28_input_sync_blk[23] | proc_28_output_sync_blk[23]);
    assign proc_28_data_FIFO_blk[24] = 1'b0;
    assign proc_28_data_PIPO_blk[24] = 1'b0;
    assign proc_28_start_FIFO_blk[24] = 1'b0;
    assign proc_28_TLF_FIFO_blk[24] = 1'b0;
    assign proc_28_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_28_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_28[24] = dl_detect_out ? proc_dep_vld_vec_28_reg[24] : (proc_28_data_FIFO_blk[24] | proc_28_data_PIPO_blk[24] | proc_28_start_FIFO_blk[24] | proc_28_TLF_FIFO_blk[24] | proc_28_input_sync_blk[24] | proc_28_output_sync_blk[24]);
    assign proc_28_data_FIFO_blk[25] = 1'b0;
    assign proc_28_data_PIPO_blk[25] = 1'b0;
    assign proc_28_start_FIFO_blk[25] = 1'b0;
    assign proc_28_TLF_FIFO_blk[25] = 1'b0;
    assign proc_28_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_28_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_28[25] = dl_detect_out ? proc_dep_vld_vec_28_reg[25] : (proc_28_data_FIFO_blk[25] | proc_28_data_PIPO_blk[25] | proc_28_start_FIFO_blk[25] | proc_28_TLF_FIFO_blk[25] | proc_28_input_sync_blk[25] | proc_28_output_sync_blk[25]);
    assign proc_28_data_FIFO_blk[26] = 1'b0;
    assign proc_28_data_PIPO_blk[26] = 1'b0;
    assign proc_28_start_FIFO_blk[26] = 1'b0;
    assign proc_28_TLF_FIFO_blk[26] = 1'b0;
    assign proc_28_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_28_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_28[26] = dl_detect_out ? proc_dep_vld_vec_28_reg[26] : (proc_28_data_FIFO_blk[26] | proc_28_data_PIPO_blk[26] | proc_28_start_FIFO_blk[26] | proc_28_TLF_FIFO_blk[26] | proc_28_input_sync_blk[26] | proc_28_output_sync_blk[26]);
    assign proc_28_data_FIFO_blk[27] = 1'b0;
    assign proc_28_data_PIPO_blk[27] = 1'b0;
    assign proc_28_start_FIFO_blk[27] = 1'b0;
    assign proc_28_TLF_FIFO_blk[27] = 1'b0;
    assign proc_28_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_28_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_28[27] = dl_detect_out ? proc_dep_vld_vec_28_reg[27] : (proc_28_data_FIFO_blk[27] | proc_28_data_PIPO_blk[27] | proc_28_start_FIFO_blk[27] | proc_28_TLF_FIFO_blk[27] | proc_28_input_sync_blk[27] | proc_28_output_sync_blk[27]);
    assign proc_28_data_FIFO_blk[28] = 1'b0;
    assign proc_28_data_PIPO_blk[28] = 1'b0;
    assign proc_28_start_FIFO_blk[28] = 1'b0;
    assign proc_28_TLF_FIFO_blk[28] = 1'b0;
    assign proc_28_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_28_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_28[28] = dl_detect_out ? proc_dep_vld_vec_28_reg[28] : (proc_28_data_FIFO_blk[28] | proc_28_data_PIPO_blk[28] | proc_28_start_FIFO_blk[28] | proc_28_TLF_FIFO_blk[28] | proc_28_input_sync_blk[28] | proc_28_output_sync_blk[28]);
    assign proc_28_data_FIFO_blk[29] = 1'b0;
    assign proc_28_data_PIPO_blk[29] = 1'b0;
    assign proc_28_start_FIFO_blk[29] = 1'b0;
    assign proc_28_TLF_FIFO_blk[29] = 1'b0;
    assign proc_28_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_28_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_28[29] = dl_detect_out ? proc_dep_vld_vec_28_reg[29] : (proc_28_data_FIFO_blk[29] | proc_28_data_PIPO_blk[29] | proc_28_start_FIFO_blk[29] | proc_28_TLF_FIFO_blk[29] | proc_28_input_sync_blk[29] | proc_28_output_sync_blk[29]);
    assign proc_28_data_FIFO_blk[30] = 1'b0;
    assign proc_28_data_PIPO_blk[30] = 1'b0;
    assign proc_28_start_FIFO_blk[30] = 1'b0;
    assign proc_28_TLF_FIFO_blk[30] = 1'b0;
    assign proc_28_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_28_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_28[30] = dl_detect_out ? proc_dep_vld_vec_28_reg[30] : (proc_28_data_FIFO_blk[30] | proc_28_data_PIPO_blk[30] | proc_28_start_FIFO_blk[30] | proc_28_TLF_FIFO_blk[30] | proc_28_input_sync_blk[30] | proc_28_output_sync_blk[30]);
    assign proc_28_data_FIFO_blk[31] = 1'b0;
    assign proc_28_data_PIPO_blk[31] = 1'b0;
    assign proc_28_start_FIFO_blk[31] = 1'b0;
    assign proc_28_TLF_FIFO_blk[31] = 1'b0;
    assign proc_28_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_28_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_28[31] = dl_detect_out ? proc_dep_vld_vec_28_reg[31] : (proc_28_data_FIFO_blk[31] | proc_28_data_PIPO_blk[31] | proc_28_start_FIFO_blk[31] | proc_28_TLF_FIFO_blk[31] | proc_28_input_sync_blk[31] | proc_28_output_sync_blk[31]);
    assign proc_28_data_FIFO_blk[32] = 1'b0;
    assign proc_28_data_PIPO_blk[32] = 1'b0;
    assign proc_28_start_FIFO_blk[32] = 1'b0;
    assign proc_28_TLF_FIFO_blk[32] = 1'b0;
    assign proc_28_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_23_U0_ap_ready & ProcessingElement_23_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_28_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_28[32] = dl_detect_out ? proc_dep_vld_vec_28_reg[32] : (proc_28_data_FIFO_blk[32] | proc_28_data_PIPO_blk[32] | proc_28_start_FIFO_blk[32] | proc_28_TLF_FIFO_blk[32] | proc_28_input_sync_blk[32] | proc_28_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_28_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_28_reg <= proc_dep_vld_vec_28;
        end
    end
    assign in_chan_dep_vld_vec_28[0] = dep_chan_vld_0_28;
    assign in_chan_dep_data_vec_28[39 : 0] = dep_chan_data_0_28;
    assign token_in_vec_28[0] = token_0_28;
    assign in_chan_dep_vld_vec_28[1] = dep_chan_vld_1_28;
    assign in_chan_dep_data_vec_28[79 : 40] = dep_chan_data_1_28;
    assign token_in_vec_28[1] = token_1_28;
    assign in_chan_dep_vld_vec_28[2] = dep_chan_vld_3_28;
    assign in_chan_dep_data_vec_28[119 : 80] = dep_chan_data_3_28;
    assign token_in_vec_28[2] = token_3_28;
    assign in_chan_dep_vld_vec_28[3] = dep_chan_vld_6_28;
    assign in_chan_dep_data_vec_28[159 : 120] = dep_chan_data_6_28;
    assign token_in_vec_28[3] = token_6_28;
    assign in_chan_dep_vld_vec_28[4] = dep_chan_vld_7_28;
    assign in_chan_dep_data_vec_28[199 : 160] = dep_chan_data_7_28;
    assign token_in_vec_28[4] = token_7_28;
    assign in_chan_dep_vld_vec_28[5] = dep_chan_vld_8_28;
    assign in_chan_dep_data_vec_28[239 : 200] = dep_chan_data_8_28;
    assign token_in_vec_28[5] = token_8_28;
    assign in_chan_dep_vld_vec_28[6] = dep_chan_vld_9_28;
    assign in_chan_dep_data_vec_28[279 : 240] = dep_chan_data_9_28;
    assign token_in_vec_28[6] = token_9_28;
    assign in_chan_dep_vld_vec_28[7] = dep_chan_vld_10_28;
    assign in_chan_dep_data_vec_28[319 : 280] = dep_chan_data_10_28;
    assign token_in_vec_28[7] = token_10_28;
    assign in_chan_dep_vld_vec_28[8] = dep_chan_vld_11_28;
    assign in_chan_dep_data_vec_28[359 : 320] = dep_chan_data_11_28;
    assign token_in_vec_28[8] = token_11_28;
    assign in_chan_dep_vld_vec_28[9] = dep_chan_vld_12_28;
    assign in_chan_dep_data_vec_28[399 : 360] = dep_chan_data_12_28;
    assign token_in_vec_28[9] = token_12_28;
    assign in_chan_dep_vld_vec_28[10] = dep_chan_vld_13_28;
    assign in_chan_dep_data_vec_28[439 : 400] = dep_chan_data_13_28;
    assign token_in_vec_28[10] = token_13_28;
    assign in_chan_dep_vld_vec_28[11] = dep_chan_vld_14_28;
    assign in_chan_dep_data_vec_28[479 : 440] = dep_chan_data_14_28;
    assign token_in_vec_28[11] = token_14_28;
    assign in_chan_dep_vld_vec_28[12] = dep_chan_vld_15_28;
    assign in_chan_dep_data_vec_28[519 : 480] = dep_chan_data_15_28;
    assign token_in_vec_28[12] = token_15_28;
    assign in_chan_dep_vld_vec_28[13] = dep_chan_vld_16_28;
    assign in_chan_dep_data_vec_28[559 : 520] = dep_chan_data_16_28;
    assign token_in_vec_28[13] = token_16_28;
    assign in_chan_dep_vld_vec_28[14] = dep_chan_vld_17_28;
    assign in_chan_dep_data_vec_28[599 : 560] = dep_chan_data_17_28;
    assign token_in_vec_28[14] = token_17_28;
    assign in_chan_dep_vld_vec_28[15] = dep_chan_vld_18_28;
    assign in_chan_dep_data_vec_28[639 : 600] = dep_chan_data_18_28;
    assign token_in_vec_28[15] = token_18_28;
    assign in_chan_dep_vld_vec_28[16] = dep_chan_vld_19_28;
    assign in_chan_dep_data_vec_28[679 : 640] = dep_chan_data_19_28;
    assign token_in_vec_28[16] = token_19_28;
    assign in_chan_dep_vld_vec_28[17] = dep_chan_vld_20_28;
    assign in_chan_dep_data_vec_28[719 : 680] = dep_chan_data_20_28;
    assign token_in_vec_28[17] = token_20_28;
    assign in_chan_dep_vld_vec_28[18] = dep_chan_vld_21_28;
    assign in_chan_dep_data_vec_28[759 : 720] = dep_chan_data_21_28;
    assign token_in_vec_28[18] = token_21_28;
    assign in_chan_dep_vld_vec_28[19] = dep_chan_vld_22_28;
    assign in_chan_dep_data_vec_28[799 : 760] = dep_chan_data_22_28;
    assign token_in_vec_28[19] = token_22_28;
    assign in_chan_dep_vld_vec_28[20] = dep_chan_vld_23_28;
    assign in_chan_dep_data_vec_28[839 : 800] = dep_chan_data_23_28;
    assign token_in_vec_28[20] = token_23_28;
    assign in_chan_dep_vld_vec_28[21] = dep_chan_vld_24_28;
    assign in_chan_dep_data_vec_28[879 : 840] = dep_chan_data_24_28;
    assign token_in_vec_28[21] = token_24_28;
    assign in_chan_dep_vld_vec_28[22] = dep_chan_vld_25_28;
    assign in_chan_dep_data_vec_28[919 : 880] = dep_chan_data_25_28;
    assign token_in_vec_28[22] = token_25_28;
    assign in_chan_dep_vld_vec_28[23] = dep_chan_vld_26_28;
    assign in_chan_dep_data_vec_28[959 : 920] = dep_chan_data_26_28;
    assign token_in_vec_28[23] = token_26_28;
    assign in_chan_dep_vld_vec_28[24] = dep_chan_vld_27_28;
    assign in_chan_dep_data_vec_28[999 : 960] = dep_chan_data_27_28;
    assign token_in_vec_28[24] = token_27_28;
    assign in_chan_dep_vld_vec_28[25] = dep_chan_vld_29_28;
    assign in_chan_dep_data_vec_28[1039 : 1000] = dep_chan_data_29_28;
    assign token_in_vec_28[25] = token_29_28;
    assign in_chan_dep_vld_vec_28[26] = dep_chan_vld_30_28;
    assign in_chan_dep_data_vec_28[1079 : 1040] = dep_chan_data_30_28;
    assign token_in_vec_28[26] = token_30_28;
    assign in_chan_dep_vld_vec_28[27] = dep_chan_vld_31_28;
    assign in_chan_dep_data_vec_28[1119 : 1080] = dep_chan_data_31_28;
    assign token_in_vec_28[27] = token_31_28;
    assign in_chan_dep_vld_vec_28[28] = dep_chan_vld_32_28;
    assign in_chan_dep_data_vec_28[1159 : 1120] = dep_chan_data_32_28;
    assign token_in_vec_28[28] = token_32_28;
    assign in_chan_dep_vld_vec_28[29] = dep_chan_vld_33_28;
    assign in_chan_dep_data_vec_28[1199 : 1160] = dep_chan_data_33_28;
    assign token_in_vec_28[29] = token_33_28;
    assign in_chan_dep_vld_vec_28[30] = dep_chan_vld_34_28;
    assign in_chan_dep_data_vec_28[1239 : 1200] = dep_chan_data_34_28;
    assign token_in_vec_28[30] = token_34_28;
    assign in_chan_dep_vld_vec_28[31] = dep_chan_vld_35_28;
    assign in_chan_dep_data_vec_28[1279 : 1240] = dep_chan_data_35_28;
    assign token_in_vec_28[31] = token_35_28;
    assign in_chan_dep_vld_vec_28[32] = dep_chan_vld_36_28;
    assign in_chan_dep_data_vec_28[1319 : 1280] = dep_chan_data_36_28;
    assign token_in_vec_28[32] = token_36_28;
    assign dep_chan_vld_28_27 = out_chan_dep_vld_vec_28[0];
    assign dep_chan_data_28_27 = out_chan_dep_data_28;
    assign token_28_27 = token_out_vec_28[0];
    assign dep_chan_vld_28_29 = out_chan_dep_vld_vec_28[1];
    assign dep_chan_data_28_29 = out_chan_dep_data_28;
    assign token_28_29 = token_out_vec_28[1];
    assign dep_chan_vld_28_0 = out_chan_dep_vld_vec_28[2];
    assign dep_chan_data_28_0 = out_chan_dep_data_28;
    assign token_28_0 = token_out_vec_28[2];
    assign dep_chan_vld_28_1 = out_chan_dep_vld_vec_28[3];
    assign dep_chan_data_28_1 = out_chan_dep_data_28;
    assign token_28_1 = token_out_vec_28[3];
    assign dep_chan_vld_28_3 = out_chan_dep_vld_vec_28[4];
    assign dep_chan_data_28_3 = out_chan_dep_data_28;
    assign token_28_3 = token_out_vec_28[4];
    assign dep_chan_vld_28_6 = out_chan_dep_vld_vec_28[5];
    assign dep_chan_data_28_6 = out_chan_dep_data_28;
    assign token_28_6 = token_out_vec_28[5];
    assign dep_chan_vld_28_7 = out_chan_dep_vld_vec_28[6];
    assign dep_chan_data_28_7 = out_chan_dep_data_28;
    assign token_28_7 = token_out_vec_28[6];
    assign dep_chan_vld_28_8 = out_chan_dep_vld_vec_28[7];
    assign dep_chan_data_28_8 = out_chan_dep_data_28;
    assign token_28_8 = token_out_vec_28[7];
    assign dep_chan_vld_28_9 = out_chan_dep_vld_vec_28[8];
    assign dep_chan_data_28_9 = out_chan_dep_data_28;
    assign token_28_9 = token_out_vec_28[8];
    assign dep_chan_vld_28_10 = out_chan_dep_vld_vec_28[9];
    assign dep_chan_data_28_10 = out_chan_dep_data_28;
    assign token_28_10 = token_out_vec_28[9];
    assign dep_chan_vld_28_11 = out_chan_dep_vld_vec_28[10];
    assign dep_chan_data_28_11 = out_chan_dep_data_28;
    assign token_28_11 = token_out_vec_28[10];
    assign dep_chan_vld_28_12 = out_chan_dep_vld_vec_28[11];
    assign dep_chan_data_28_12 = out_chan_dep_data_28;
    assign token_28_12 = token_out_vec_28[11];
    assign dep_chan_vld_28_13 = out_chan_dep_vld_vec_28[12];
    assign dep_chan_data_28_13 = out_chan_dep_data_28;
    assign token_28_13 = token_out_vec_28[12];
    assign dep_chan_vld_28_14 = out_chan_dep_vld_vec_28[13];
    assign dep_chan_data_28_14 = out_chan_dep_data_28;
    assign token_28_14 = token_out_vec_28[13];
    assign dep_chan_vld_28_15 = out_chan_dep_vld_vec_28[14];
    assign dep_chan_data_28_15 = out_chan_dep_data_28;
    assign token_28_15 = token_out_vec_28[14];
    assign dep_chan_vld_28_16 = out_chan_dep_vld_vec_28[15];
    assign dep_chan_data_28_16 = out_chan_dep_data_28;
    assign token_28_16 = token_out_vec_28[15];
    assign dep_chan_vld_28_17 = out_chan_dep_vld_vec_28[16];
    assign dep_chan_data_28_17 = out_chan_dep_data_28;
    assign token_28_17 = token_out_vec_28[16];
    assign dep_chan_vld_28_18 = out_chan_dep_vld_vec_28[17];
    assign dep_chan_data_28_18 = out_chan_dep_data_28;
    assign token_28_18 = token_out_vec_28[17];
    assign dep_chan_vld_28_19 = out_chan_dep_vld_vec_28[18];
    assign dep_chan_data_28_19 = out_chan_dep_data_28;
    assign token_28_19 = token_out_vec_28[18];
    assign dep_chan_vld_28_20 = out_chan_dep_vld_vec_28[19];
    assign dep_chan_data_28_20 = out_chan_dep_data_28;
    assign token_28_20 = token_out_vec_28[19];
    assign dep_chan_vld_28_21 = out_chan_dep_vld_vec_28[20];
    assign dep_chan_data_28_21 = out_chan_dep_data_28;
    assign token_28_21 = token_out_vec_28[20];
    assign dep_chan_vld_28_22 = out_chan_dep_vld_vec_28[21];
    assign dep_chan_data_28_22 = out_chan_dep_data_28;
    assign token_28_22 = token_out_vec_28[21];
    assign dep_chan_vld_28_23 = out_chan_dep_vld_vec_28[22];
    assign dep_chan_data_28_23 = out_chan_dep_data_28;
    assign token_28_23 = token_out_vec_28[22];
    assign dep_chan_vld_28_24 = out_chan_dep_vld_vec_28[23];
    assign dep_chan_data_28_24 = out_chan_dep_data_28;
    assign token_28_24 = token_out_vec_28[23];
    assign dep_chan_vld_28_25 = out_chan_dep_vld_vec_28[24];
    assign dep_chan_data_28_25 = out_chan_dep_data_28;
    assign token_28_25 = token_out_vec_28[24];
    assign dep_chan_vld_28_26 = out_chan_dep_vld_vec_28[25];
    assign dep_chan_data_28_26 = out_chan_dep_data_28;
    assign token_28_26 = token_out_vec_28[25];
    assign dep_chan_vld_28_30 = out_chan_dep_vld_vec_28[26];
    assign dep_chan_data_28_30 = out_chan_dep_data_28;
    assign token_28_30 = token_out_vec_28[26];
    assign dep_chan_vld_28_31 = out_chan_dep_vld_vec_28[27];
    assign dep_chan_data_28_31 = out_chan_dep_data_28;
    assign token_28_31 = token_out_vec_28[27];
    assign dep_chan_vld_28_32 = out_chan_dep_vld_vec_28[28];
    assign dep_chan_data_28_32 = out_chan_dep_data_28;
    assign token_28_32 = token_out_vec_28[28];
    assign dep_chan_vld_28_33 = out_chan_dep_vld_vec_28[29];
    assign dep_chan_data_28_33 = out_chan_dep_data_28;
    assign token_28_33 = token_out_vec_28[29];
    assign dep_chan_vld_28_34 = out_chan_dep_vld_vec_28[30];
    assign dep_chan_data_28_34 = out_chan_dep_data_28;
    assign token_28_34 = token_out_vec_28[30];
    assign dep_chan_vld_28_35 = out_chan_dep_vld_vec_28[31];
    assign dep_chan_data_28_35 = out_chan_dep_data_28;
    assign token_28_35 = token_out_vec_28[31];
    assign dep_chan_vld_28_36 = out_chan_dep_vld_vec_28[32];
    assign dep_chan_data_28_36 = out_chan_dep_data_28;
    assign token_28_36 = token_out_vec_28[32];

    // Process: ProcessingElement_24_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 29, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_29 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_29),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_29),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_29),
        .token_in_vec(token_in_vec_29),
        .dl_detect_in(dl_detect_out),
        .origin(origin[29]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_29),
        .out_chan_dep_data(out_chan_dep_data_29),
        .token_out_vec(token_out_vec_29),
        .dl_detect_out(dl_in_vec[29]));

    assign proc_29_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_23_blk_n) | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_23_blk_n) | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_WriteC_Flattened_fu_179.cPipes_23_blk_n);
    assign proc_29_data_PIPO_blk[0] = 1'b0;
    assign proc_29_start_FIFO_blk[0] = 1'b0;
    assign proc_29_TLF_FIFO_blk[0] = 1'b0;
    assign proc_29_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_29_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_29[0] = dl_detect_out ? proc_dep_vld_vec_29_reg[0] : (proc_29_data_FIFO_blk[0] | proc_29_data_PIPO_blk[0] | proc_29_start_FIFO_blk[0] | proc_29_TLF_FIFO_blk[0] | proc_29_input_sync_blk[0] | proc_29_output_sync_blk[0]);
    assign proc_29_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_24_blk_n) | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_24_blk_n) | (~ProcessingElement_24_U0.grp_ProcessingElement_24_Pipeline_WriteC_Flattened_fu_179.cPipes_24_blk_n);
    assign proc_29_data_PIPO_blk[1] = 1'b0;
    assign proc_29_start_FIFO_blk[1] = 1'b0;
    assign proc_29_TLF_FIFO_blk[1] = 1'b0;
    assign proc_29_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_29_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_29[1] = dl_detect_out ? proc_dep_vld_vec_29_reg[1] : (proc_29_data_FIFO_blk[1] | proc_29_data_PIPO_blk[1] | proc_29_start_FIFO_blk[1] | proc_29_TLF_FIFO_blk[1] | proc_29_input_sync_blk[1] | proc_29_output_sync_blk[1]);
    assign proc_29_data_FIFO_blk[2] = 1'b0;
    assign proc_29_data_PIPO_blk[2] = 1'b0;
    assign proc_29_start_FIFO_blk[2] = 1'b0;
    assign proc_29_TLF_FIFO_blk[2] = 1'b0;
    assign proc_29_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_29_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_29[2] = dl_detect_out ? proc_dep_vld_vec_29_reg[2] : (proc_29_data_FIFO_blk[2] | proc_29_data_PIPO_blk[2] | proc_29_start_FIFO_blk[2] | proc_29_TLF_FIFO_blk[2] | proc_29_input_sync_blk[2] | proc_29_output_sync_blk[2]);
    assign proc_29_data_FIFO_blk[3] = 1'b0;
    assign proc_29_data_PIPO_blk[3] = 1'b0;
    assign proc_29_start_FIFO_blk[3] = 1'b0;
    assign proc_29_TLF_FIFO_blk[3] = 1'b0;
    assign proc_29_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_29_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_29[3] = dl_detect_out ? proc_dep_vld_vec_29_reg[3] : (proc_29_data_FIFO_blk[3] | proc_29_data_PIPO_blk[3] | proc_29_start_FIFO_blk[3] | proc_29_TLF_FIFO_blk[3] | proc_29_input_sync_blk[3] | proc_29_output_sync_blk[3]);
    assign proc_29_data_FIFO_blk[4] = 1'b0;
    assign proc_29_data_PIPO_blk[4] = 1'b0;
    assign proc_29_start_FIFO_blk[4] = 1'b0;
    assign proc_29_TLF_FIFO_blk[4] = 1'b0;
    assign proc_29_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_29_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_29[4] = dl_detect_out ? proc_dep_vld_vec_29_reg[4] : (proc_29_data_FIFO_blk[4] | proc_29_data_PIPO_blk[4] | proc_29_start_FIFO_blk[4] | proc_29_TLF_FIFO_blk[4] | proc_29_input_sync_blk[4] | proc_29_output_sync_blk[4]);
    assign proc_29_data_FIFO_blk[5] = 1'b0;
    assign proc_29_data_PIPO_blk[5] = 1'b0;
    assign proc_29_start_FIFO_blk[5] = 1'b0;
    assign proc_29_TLF_FIFO_blk[5] = 1'b0;
    assign proc_29_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_29_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_29[5] = dl_detect_out ? proc_dep_vld_vec_29_reg[5] : (proc_29_data_FIFO_blk[5] | proc_29_data_PIPO_blk[5] | proc_29_start_FIFO_blk[5] | proc_29_TLF_FIFO_blk[5] | proc_29_input_sync_blk[5] | proc_29_output_sync_blk[5]);
    assign proc_29_data_FIFO_blk[6] = 1'b0;
    assign proc_29_data_PIPO_blk[6] = 1'b0;
    assign proc_29_start_FIFO_blk[6] = 1'b0;
    assign proc_29_TLF_FIFO_blk[6] = 1'b0;
    assign proc_29_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_29_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_29[6] = dl_detect_out ? proc_dep_vld_vec_29_reg[6] : (proc_29_data_FIFO_blk[6] | proc_29_data_PIPO_blk[6] | proc_29_start_FIFO_blk[6] | proc_29_TLF_FIFO_blk[6] | proc_29_input_sync_blk[6] | proc_29_output_sync_blk[6]);
    assign proc_29_data_FIFO_blk[7] = 1'b0;
    assign proc_29_data_PIPO_blk[7] = 1'b0;
    assign proc_29_start_FIFO_blk[7] = 1'b0;
    assign proc_29_TLF_FIFO_blk[7] = 1'b0;
    assign proc_29_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_29_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_29[7] = dl_detect_out ? proc_dep_vld_vec_29_reg[7] : (proc_29_data_FIFO_blk[7] | proc_29_data_PIPO_blk[7] | proc_29_start_FIFO_blk[7] | proc_29_TLF_FIFO_blk[7] | proc_29_input_sync_blk[7] | proc_29_output_sync_blk[7]);
    assign proc_29_data_FIFO_blk[8] = 1'b0;
    assign proc_29_data_PIPO_blk[8] = 1'b0;
    assign proc_29_start_FIFO_blk[8] = 1'b0;
    assign proc_29_TLF_FIFO_blk[8] = 1'b0;
    assign proc_29_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_29_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_29[8] = dl_detect_out ? proc_dep_vld_vec_29_reg[8] : (proc_29_data_FIFO_blk[8] | proc_29_data_PIPO_blk[8] | proc_29_start_FIFO_blk[8] | proc_29_TLF_FIFO_blk[8] | proc_29_input_sync_blk[8] | proc_29_output_sync_blk[8]);
    assign proc_29_data_FIFO_blk[9] = 1'b0;
    assign proc_29_data_PIPO_blk[9] = 1'b0;
    assign proc_29_start_FIFO_blk[9] = 1'b0;
    assign proc_29_TLF_FIFO_blk[9] = 1'b0;
    assign proc_29_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_29_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_29[9] = dl_detect_out ? proc_dep_vld_vec_29_reg[9] : (proc_29_data_FIFO_blk[9] | proc_29_data_PIPO_blk[9] | proc_29_start_FIFO_blk[9] | proc_29_TLF_FIFO_blk[9] | proc_29_input_sync_blk[9] | proc_29_output_sync_blk[9]);
    assign proc_29_data_FIFO_blk[10] = 1'b0;
    assign proc_29_data_PIPO_blk[10] = 1'b0;
    assign proc_29_start_FIFO_blk[10] = 1'b0;
    assign proc_29_TLF_FIFO_blk[10] = 1'b0;
    assign proc_29_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_29_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_29[10] = dl_detect_out ? proc_dep_vld_vec_29_reg[10] : (proc_29_data_FIFO_blk[10] | proc_29_data_PIPO_blk[10] | proc_29_start_FIFO_blk[10] | proc_29_TLF_FIFO_blk[10] | proc_29_input_sync_blk[10] | proc_29_output_sync_blk[10]);
    assign proc_29_data_FIFO_blk[11] = 1'b0;
    assign proc_29_data_PIPO_blk[11] = 1'b0;
    assign proc_29_start_FIFO_blk[11] = 1'b0;
    assign proc_29_TLF_FIFO_blk[11] = 1'b0;
    assign proc_29_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_29_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_29[11] = dl_detect_out ? proc_dep_vld_vec_29_reg[11] : (proc_29_data_FIFO_blk[11] | proc_29_data_PIPO_blk[11] | proc_29_start_FIFO_blk[11] | proc_29_TLF_FIFO_blk[11] | proc_29_input_sync_blk[11] | proc_29_output_sync_blk[11]);
    assign proc_29_data_FIFO_blk[12] = 1'b0;
    assign proc_29_data_PIPO_blk[12] = 1'b0;
    assign proc_29_start_FIFO_blk[12] = 1'b0;
    assign proc_29_TLF_FIFO_blk[12] = 1'b0;
    assign proc_29_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_29_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_29[12] = dl_detect_out ? proc_dep_vld_vec_29_reg[12] : (proc_29_data_FIFO_blk[12] | proc_29_data_PIPO_blk[12] | proc_29_start_FIFO_blk[12] | proc_29_TLF_FIFO_blk[12] | proc_29_input_sync_blk[12] | proc_29_output_sync_blk[12]);
    assign proc_29_data_FIFO_blk[13] = 1'b0;
    assign proc_29_data_PIPO_blk[13] = 1'b0;
    assign proc_29_start_FIFO_blk[13] = 1'b0;
    assign proc_29_TLF_FIFO_blk[13] = 1'b0;
    assign proc_29_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_29_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_29[13] = dl_detect_out ? proc_dep_vld_vec_29_reg[13] : (proc_29_data_FIFO_blk[13] | proc_29_data_PIPO_blk[13] | proc_29_start_FIFO_blk[13] | proc_29_TLF_FIFO_blk[13] | proc_29_input_sync_blk[13] | proc_29_output_sync_blk[13]);
    assign proc_29_data_FIFO_blk[14] = 1'b0;
    assign proc_29_data_PIPO_blk[14] = 1'b0;
    assign proc_29_start_FIFO_blk[14] = 1'b0;
    assign proc_29_TLF_FIFO_blk[14] = 1'b0;
    assign proc_29_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_29_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_29[14] = dl_detect_out ? proc_dep_vld_vec_29_reg[14] : (proc_29_data_FIFO_blk[14] | proc_29_data_PIPO_blk[14] | proc_29_start_FIFO_blk[14] | proc_29_TLF_FIFO_blk[14] | proc_29_input_sync_blk[14] | proc_29_output_sync_blk[14]);
    assign proc_29_data_FIFO_blk[15] = 1'b0;
    assign proc_29_data_PIPO_blk[15] = 1'b0;
    assign proc_29_start_FIFO_blk[15] = 1'b0;
    assign proc_29_TLF_FIFO_blk[15] = 1'b0;
    assign proc_29_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_29_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_29[15] = dl_detect_out ? proc_dep_vld_vec_29_reg[15] : (proc_29_data_FIFO_blk[15] | proc_29_data_PIPO_blk[15] | proc_29_start_FIFO_blk[15] | proc_29_TLF_FIFO_blk[15] | proc_29_input_sync_blk[15] | proc_29_output_sync_blk[15]);
    assign proc_29_data_FIFO_blk[16] = 1'b0;
    assign proc_29_data_PIPO_blk[16] = 1'b0;
    assign proc_29_start_FIFO_blk[16] = 1'b0;
    assign proc_29_TLF_FIFO_blk[16] = 1'b0;
    assign proc_29_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_29_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_29[16] = dl_detect_out ? proc_dep_vld_vec_29_reg[16] : (proc_29_data_FIFO_blk[16] | proc_29_data_PIPO_blk[16] | proc_29_start_FIFO_blk[16] | proc_29_TLF_FIFO_blk[16] | proc_29_input_sync_blk[16] | proc_29_output_sync_blk[16]);
    assign proc_29_data_FIFO_blk[17] = 1'b0;
    assign proc_29_data_PIPO_blk[17] = 1'b0;
    assign proc_29_start_FIFO_blk[17] = 1'b0;
    assign proc_29_TLF_FIFO_blk[17] = 1'b0;
    assign proc_29_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_29_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_29[17] = dl_detect_out ? proc_dep_vld_vec_29_reg[17] : (proc_29_data_FIFO_blk[17] | proc_29_data_PIPO_blk[17] | proc_29_start_FIFO_blk[17] | proc_29_TLF_FIFO_blk[17] | proc_29_input_sync_blk[17] | proc_29_output_sync_blk[17]);
    assign proc_29_data_FIFO_blk[18] = 1'b0;
    assign proc_29_data_PIPO_blk[18] = 1'b0;
    assign proc_29_start_FIFO_blk[18] = 1'b0;
    assign proc_29_TLF_FIFO_blk[18] = 1'b0;
    assign proc_29_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_29_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_29[18] = dl_detect_out ? proc_dep_vld_vec_29_reg[18] : (proc_29_data_FIFO_blk[18] | proc_29_data_PIPO_blk[18] | proc_29_start_FIFO_blk[18] | proc_29_TLF_FIFO_blk[18] | proc_29_input_sync_blk[18] | proc_29_output_sync_blk[18]);
    assign proc_29_data_FIFO_blk[19] = 1'b0;
    assign proc_29_data_PIPO_blk[19] = 1'b0;
    assign proc_29_start_FIFO_blk[19] = 1'b0;
    assign proc_29_TLF_FIFO_blk[19] = 1'b0;
    assign proc_29_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_29_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_29[19] = dl_detect_out ? proc_dep_vld_vec_29_reg[19] : (proc_29_data_FIFO_blk[19] | proc_29_data_PIPO_blk[19] | proc_29_start_FIFO_blk[19] | proc_29_TLF_FIFO_blk[19] | proc_29_input_sync_blk[19] | proc_29_output_sync_blk[19]);
    assign proc_29_data_FIFO_blk[20] = 1'b0;
    assign proc_29_data_PIPO_blk[20] = 1'b0;
    assign proc_29_start_FIFO_blk[20] = 1'b0;
    assign proc_29_TLF_FIFO_blk[20] = 1'b0;
    assign proc_29_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_29_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_29[20] = dl_detect_out ? proc_dep_vld_vec_29_reg[20] : (proc_29_data_FIFO_blk[20] | proc_29_data_PIPO_blk[20] | proc_29_start_FIFO_blk[20] | proc_29_TLF_FIFO_blk[20] | proc_29_input_sync_blk[20] | proc_29_output_sync_blk[20]);
    assign proc_29_data_FIFO_blk[21] = 1'b0;
    assign proc_29_data_PIPO_blk[21] = 1'b0;
    assign proc_29_start_FIFO_blk[21] = 1'b0;
    assign proc_29_TLF_FIFO_blk[21] = 1'b0;
    assign proc_29_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_29_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_29[21] = dl_detect_out ? proc_dep_vld_vec_29_reg[21] : (proc_29_data_FIFO_blk[21] | proc_29_data_PIPO_blk[21] | proc_29_start_FIFO_blk[21] | proc_29_TLF_FIFO_blk[21] | proc_29_input_sync_blk[21] | proc_29_output_sync_blk[21]);
    assign proc_29_data_FIFO_blk[22] = 1'b0;
    assign proc_29_data_PIPO_blk[22] = 1'b0;
    assign proc_29_start_FIFO_blk[22] = 1'b0;
    assign proc_29_TLF_FIFO_blk[22] = 1'b0;
    assign proc_29_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_29_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_29[22] = dl_detect_out ? proc_dep_vld_vec_29_reg[22] : (proc_29_data_FIFO_blk[22] | proc_29_data_PIPO_blk[22] | proc_29_start_FIFO_blk[22] | proc_29_TLF_FIFO_blk[22] | proc_29_input_sync_blk[22] | proc_29_output_sync_blk[22]);
    assign proc_29_data_FIFO_blk[23] = 1'b0;
    assign proc_29_data_PIPO_blk[23] = 1'b0;
    assign proc_29_start_FIFO_blk[23] = 1'b0;
    assign proc_29_TLF_FIFO_blk[23] = 1'b0;
    assign proc_29_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_29_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_29[23] = dl_detect_out ? proc_dep_vld_vec_29_reg[23] : (proc_29_data_FIFO_blk[23] | proc_29_data_PIPO_blk[23] | proc_29_start_FIFO_blk[23] | proc_29_TLF_FIFO_blk[23] | proc_29_input_sync_blk[23] | proc_29_output_sync_blk[23]);
    assign proc_29_data_FIFO_blk[24] = 1'b0;
    assign proc_29_data_PIPO_blk[24] = 1'b0;
    assign proc_29_start_FIFO_blk[24] = 1'b0;
    assign proc_29_TLF_FIFO_blk[24] = 1'b0;
    assign proc_29_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_29_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_29[24] = dl_detect_out ? proc_dep_vld_vec_29_reg[24] : (proc_29_data_FIFO_blk[24] | proc_29_data_PIPO_blk[24] | proc_29_start_FIFO_blk[24] | proc_29_TLF_FIFO_blk[24] | proc_29_input_sync_blk[24] | proc_29_output_sync_blk[24]);
    assign proc_29_data_FIFO_blk[25] = 1'b0;
    assign proc_29_data_PIPO_blk[25] = 1'b0;
    assign proc_29_start_FIFO_blk[25] = 1'b0;
    assign proc_29_TLF_FIFO_blk[25] = 1'b0;
    assign proc_29_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_29_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_29[25] = dl_detect_out ? proc_dep_vld_vec_29_reg[25] : (proc_29_data_FIFO_blk[25] | proc_29_data_PIPO_blk[25] | proc_29_start_FIFO_blk[25] | proc_29_TLF_FIFO_blk[25] | proc_29_input_sync_blk[25] | proc_29_output_sync_blk[25]);
    assign proc_29_data_FIFO_blk[26] = 1'b0;
    assign proc_29_data_PIPO_blk[26] = 1'b0;
    assign proc_29_start_FIFO_blk[26] = 1'b0;
    assign proc_29_TLF_FIFO_blk[26] = 1'b0;
    assign proc_29_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_29_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_29[26] = dl_detect_out ? proc_dep_vld_vec_29_reg[26] : (proc_29_data_FIFO_blk[26] | proc_29_data_PIPO_blk[26] | proc_29_start_FIFO_blk[26] | proc_29_TLF_FIFO_blk[26] | proc_29_input_sync_blk[26] | proc_29_output_sync_blk[26]);
    assign proc_29_data_FIFO_blk[27] = 1'b0;
    assign proc_29_data_PIPO_blk[27] = 1'b0;
    assign proc_29_start_FIFO_blk[27] = 1'b0;
    assign proc_29_TLF_FIFO_blk[27] = 1'b0;
    assign proc_29_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_29_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_29[27] = dl_detect_out ? proc_dep_vld_vec_29_reg[27] : (proc_29_data_FIFO_blk[27] | proc_29_data_PIPO_blk[27] | proc_29_start_FIFO_blk[27] | proc_29_TLF_FIFO_blk[27] | proc_29_input_sync_blk[27] | proc_29_output_sync_blk[27]);
    assign proc_29_data_FIFO_blk[28] = 1'b0;
    assign proc_29_data_PIPO_blk[28] = 1'b0;
    assign proc_29_start_FIFO_blk[28] = 1'b0;
    assign proc_29_TLF_FIFO_blk[28] = 1'b0;
    assign proc_29_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_29_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_29[28] = dl_detect_out ? proc_dep_vld_vec_29_reg[28] : (proc_29_data_FIFO_blk[28] | proc_29_data_PIPO_blk[28] | proc_29_start_FIFO_blk[28] | proc_29_TLF_FIFO_blk[28] | proc_29_input_sync_blk[28] | proc_29_output_sync_blk[28]);
    assign proc_29_data_FIFO_blk[29] = 1'b0;
    assign proc_29_data_PIPO_blk[29] = 1'b0;
    assign proc_29_start_FIFO_blk[29] = 1'b0;
    assign proc_29_TLF_FIFO_blk[29] = 1'b0;
    assign proc_29_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_29_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_29[29] = dl_detect_out ? proc_dep_vld_vec_29_reg[29] : (proc_29_data_FIFO_blk[29] | proc_29_data_PIPO_blk[29] | proc_29_start_FIFO_blk[29] | proc_29_TLF_FIFO_blk[29] | proc_29_input_sync_blk[29] | proc_29_output_sync_blk[29]);
    assign proc_29_data_FIFO_blk[30] = 1'b0;
    assign proc_29_data_PIPO_blk[30] = 1'b0;
    assign proc_29_start_FIFO_blk[30] = 1'b0;
    assign proc_29_TLF_FIFO_blk[30] = 1'b0;
    assign proc_29_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_29_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_29[30] = dl_detect_out ? proc_dep_vld_vec_29_reg[30] : (proc_29_data_FIFO_blk[30] | proc_29_data_PIPO_blk[30] | proc_29_start_FIFO_blk[30] | proc_29_TLF_FIFO_blk[30] | proc_29_input_sync_blk[30] | proc_29_output_sync_blk[30]);
    assign proc_29_data_FIFO_blk[31] = 1'b0;
    assign proc_29_data_PIPO_blk[31] = 1'b0;
    assign proc_29_start_FIFO_blk[31] = 1'b0;
    assign proc_29_TLF_FIFO_blk[31] = 1'b0;
    assign proc_29_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_29_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_29[31] = dl_detect_out ? proc_dep_vld_vec_29_reg[31] : (proc_29_data_FIFO_blk[31] | proc_29_data_PIPO_blk[31] | proc_29_start_FIFO_blk[31] | proc_29_TLF_FIFO_blk[31] | proc_29_input_sync_blk[31] | proc_29_output_sync_blk[31]);
    assign proc_29_data_FIFO_blk[32] = 1'b0;
    assign proc_29_data_PIPO_blk[32] = 1'b0;
    assign proc_29_start_FIFO_blk[32] = 1'b0;
    assign proc_29_TLF_FIFO_blk[32] = 1'b0;
    assign proc_29_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_24_U0_ap_ready & ProcessingElement_24_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_29_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_29[32] = dl_detect_out ? proc_dep_vld_vec_29_reg[32] : (proc_29_data_FIFO_blk[32] | proc_29_data_PIPO_blk[32] | proc_29_start_FIFO_blk[32] | proc_29_TLF_FIFO_blk[32] | proc_29_input_sync_blk[32] | proc_29_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_29_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_29_reg <= proc_dep_vld_vec_29;
        end
    end
    assign in_chan_dep_vld_vec_29[0] = dep_chan_vld_0_29;
    assign in_chan_dep_data_vec_29[39 : 0] = dep_chan_data_0_29;
    assign token_in_vec_29[0] = token_0_29;
    assign in_chan_dep_vld_vec_29[1] = dep_chan_vld_1_29;
    assign in_chan_dep_data_vec_29[79 : 40] = dep_chan_data_1_29;
    assign token_in_vec_29[1] = token_1_29;
    assign in_chan_dep_vld_vec_29[2] = dep_chan_vld_3_29;
    assign in_chan_dep_data_vec_29[119 : 80] = dep_chan_data_3_29;
    assign token_in_vec_29[2] = token_3_29;
    assign in_chan_dep_vld_vec_29[3] = dep_chan_vld_6_29;
    assign in_chan_dep_data_vec_29[159 : 120] = dep_chan_data_6_29;
    assign token_in_vec_29[3] = token_6_29;
    assign in_chan_dep_vld_vec_29[4] = dep_chan_vld_7_29;
    assign in_chan_dep_data_vec_29[199 : 160] = dep_chan_data_7_29;
    assign token_in_vec_29[4] = token_7_29;
    assign in_chan_dep_vld_vec_29[5] = dep_chan_vld_8_29;
    assign in_chan_dep_data_vec_29[239 : 200] = dep_chan_data_8_29;
    assign token_in_vec_29[5] = token_8_29;
    assign in_chan_dep_vld_vec_29[6] = dep_chan_vld_9_29;
    assign in_chan_dep_data_vec_29[279 : 240] = dep_chan_data_9_29;
    assign token_in_vec_29[6] = token_9_29;
    assign in_chan_dep_vld_vec_29[7] = dep_chan_vld_10_29;
    assign in_chan_dep_data_vec_29[319 : 280] = dep_chan_data_10_29;
    assign token_in_vec_29[7] = token_10_29;
    assign in_chan_dep_vld_vec_29[8] = dep_chan_vld_11_29;
    assign in_chan_dep_data_vec_29[359 : 320] = dep_chan_data_11_29;
    assign token_in_vec_29[8] = token_11_29;
    assign in_chan_dep_vld_vec_29[9] = dep_chan_vld_12_29;
    assign in_chan_dep_data_vec_29[399 : 360] = dep_chan_data_12_29;
    assign token_in_vec_29[9] = token_12_29;
    assign in_chan_dep_vld_vec_29[10] = dep_chan_vld_13_29;
    assign in_chan_dep_data_vec_29[439 : 400] = dep_chan_data_13_29;
    assign token_in_vec_29[10] = token_13_29;
    assign in_chan_dep_vld_vec_29[11] = dep_chan_vld_14_29;
    assign in_chan_dep_data_vec_29[479 : 440] = dep_chan_data_14_29;
    assign token_in_vec_29[11] = token_14_29;
    assign in_chan_dep_vld_vec_29[12] = dep_chan_vld_15_29;
    assign in_chan_dep_data_vec_29[519 : 480] = dep_chan_data_15_29;
    assign token_in_vec_29[12] = token_15_29;
    assign in_chan_dep_vld_vec_29[13] = dep_chan_vld_16_29;
    assign in_chan_dep_data_vec_29[559 : 520] = dep_chan_data_16_29;
    assign token_in_vec_29[13] = token_16_29;
    assign in_chan_dep_vld_vec_29[14] = dep_chan_vld_17_29;
    assign in_chan_dep_data_vec_29[599 : 560] = dep_chan_data_17_29;
    assign token_in_vec_29[14] = token_17_29;
    assign in_chan_dep_vld_vec_29[15] = dep_chan_vld_18_29;
    assign in_chan_dep_data_vec_29[639 : 600] = dep_chan_data_18_29;
    assign token_in_vec_29[15] = token_18_29;
    assign in_chan_dep_vld_vec_29[16] = dep_chan_vld_19_29;
    assign in_chan_dep_data_vec_29[679 : 640] = dep_chan_data_19_29;
    assign token_in_vec_29[16] = token_19_29;
    assign in_chan_dep_vld_vec_29[17] = dep_chan_vld_20_29;
    assign in_chan_dep_data_vec_29[719 : 680] = dep_chan_data_20_29;
    assign token_in_vec_29[17] = token_20_29;
    assign in_chan_dep_vld_vec_29[18] = dep_chan_vld_21_29;
    assign in_chan_dep_data_vec_29[759 : 720] = dep_chan_data_21_29;
    assign token_in_vec_29[18] = token_21_29;
    assign in_chan_dep_vld_vec_29[19] = dep_chan_vld_22_29;
    assign in_chan_dep_data_vec_29[799 : 760] = dep_chan_data_22_29;
    assign token_in_vec_29[19] = token_22_29;
    assign in_chan_dep_vld_vec_29[20] = dep_chan_vld_23_29;
    assign in_chan_dep_data_vec_29[839 : 800] = dep_chan_data_23_29;
    assign token_in_vec_29[20] = token_23_29;
    assign in_chan_dep_vld_vec_29[21] = dep_chan_vld_24_29;
    assign in_chan_dep_data_vec_29[879 : 840] = dep_chan_data_24_29;
    assign token_in_vec_29[21] = token_24_29;
    assign in_chan_dep_vld_vec_29[22] = dep_chan_vld_25_29;
    assign in_chan_dep_data_vec_29[919 : 880] = dep_chan_data_25_29;
    assign token_in_vec_29[22] = token_25_29;
    assign in_chan_dep_vld_vec_29[23] = dep_chan_vld_26_29;
    assign in_chan_dep_data_vec_29[959 : 920] = dep_chan_data_26_29;
    assign token_in_vec_29[23] = token_26_29;
    assign in_chan_dep_vld_vec_29[24] = dep_chan_vld_27_29;
    assign in_chan_dep_data_vec_29[999 : 960] = dep_chan_data_27_29;
    assign token_in_vec_29[24] = token_27_29;
    assign in_chan_dep_vld_vec_29[25] = dep_chan_vld_28_29;
    assign in_chan_dep_data_vec_29[1039 : 1000] = dep_chan_data_28_29;
    assign token_in_vec_29[25] = token_28_29;
    assign in_chan_dep_vld_vec_29[26] = dep_chan_vld_30_29;
    assign in_chan_dep_data_vec_29[1079 : 1040] = dep_chan_data_30_29;
    assign token_in_vec_29[26] = token_30_29;
    assign in_chan_dep_vld_vec_29[27] = dep_chan_vld_31_29;
    assign in_chan_dep_data_vec_29[1119 : 1080] = dep_chan_data_31_29;
    assign token_in_vec_29[27] = token_31_29;
    assign in_chan_dep_vld_vec_29[28] = dep_chan_vld_32_29;
    assign in_chan_dep_data_vec_29[1159 : 1120] = dep_chan_data_32_29;
    assign token_in_vec_29[28] = token_32_29;
    assign in_chan_dep_vld_vec_29[29] = dep_chan_vld_33_29;
    assign in_chan_dep_data_vec_29[1199 : 1160] = dep_chan_data_33_29;
    assign token_in_vec_29[29] = token_33_29;
    assign in_chan_dep_vld_vec_29[30] = dep_chan_vld_34_29;
    assign in_chan_dep_data_vec_29[1239 : 1200] = dep_chan_data_34_29;
    assign token_in_vec_29[30] = token_34_29;
    assign in_chan_dep_vld_vec_29[31] = dep_chan_vld_35_29;
    assign in_chan_dep_data_vec_29[1279 : 1240] = dep_chan_data_35_29;
    assign token_in_vec_29[31] = token_35_29;
    assign in_chan_dep_vld_vec_29[32] = dep_chan_vld_36_29;
    assign in_chan_dep_data_vec_29[1319 : 1280] = dep_chan_data_36_29;
    assign token_in_vec_29[32] = token_36_29;
    assign dep_chan_vld_29_28 = out_chan_dep_vld_vec_29[0];
    assign dep_chan_data_29_28 = out_chan_dep_data_29;
    assign token_29_28 = token_out_vec_29[0];
    assign dep_chan_vld_29_30 = out_chan_dep_vld_vec_29[1];
    assign dep_chan_data_29_30 = out_chan_dep_data_29;
    assign token_29_30 = token_out_vec_29[1];
    assign dep_chan_vld_29_0 = out_chan_dep_vld_vec_29[2];
    assign dep_chan_data_29_0 = out_chan_dep_data_29;
    assign token_29_0 = token_out_vec_29[2];
    assign dep_chan_vld_29_1 = out_chan_dep_vld_vec_29[3];
    assign dep_chan_data_29_1 = out_chan_dep_data_29;
    assign token_29_1 = token_out_vec_29[3];
    assign dep_chan_vld_29_3 = out_chan_dep_vld_vec_29[4];
    assign dep_chan_data_29_3 = out_chan_dep_data_29;
    assign token_29_3 = token_out_vec_29[4];
    assign dep_chan_vld_29_6 = out_chan_dep_vld_vec_29[5];
    assign dep_chan_data_29_6 = out_chan_dep_data_29;
    assign token_29_6 = token_out_vec_29[5];
    assign dep_chan_vld_29_7 = out_chan_dep_vld_vec_29[6];
    assign dep_chan_data_29_7 = out_chan_dep_data_29;
    assign token_29_7 = token_out_vec_29[6];
    assign dep_chan_vld_29_8 = out_chan_dep_vld_vec_29[7];
    assign dep_chan_data_29_8 = out_chan_dep_data_29;
    assign token_29_8 = token_out_vec_29[7];
    assign dep_chan_vld_29_9 = out_chan_dep_vld_vec_29[8];
    assign dep_chan_data_29_9 = out_chan_dep_data_29;
    assign token_29_9 = token_out_vec_29[8];
    assign dep_chan_vld_29_10 = out_chan_dep_vld_vec_29[9];
    assign dep_chan_data_29_10 = out_chan_dep_data_29;
    assign token_29_10 = token_out_vec_29[9];
    assign dep_chan_vld_29_11 = out_chan_dep_vld_vec_29[10];
    assign dep_chan_data_29_11 = out_chan_dep_data_29;
    assign token_29_11 = token_out_vec_29[10];
    assign dep_chan_vld_29_12 = out_chan_dep_vld_vec_29[11];
    assign dep_chan_data_29_12 = out_chan_dep_data_29;
    assign token_29_12 = token_out_vec_29[11];
    assign dep_chan_vld_29_13 = out_chan_dep_vld_vec_29[12];
    assign dep_chan_data_29_13 = out_chan_dep_data_29;
    assign token_29_13 = token_out_vec_29[12];
    assign dep_chan_vld_29_14 = out_chan_dep_vld_vec_29[13];
    assign dep_chan_data_29_14 = out_chan_dep_data_29;
    assign token_29_14 = token_out_vec_29[13];
    assign dep_chan_vld_29_15 = out_chan_dep_vld_vec_29[14];
    assign dep_chan_data_29_15 = out_chan_dep_data_29;
    assign token_29_15 = token_out_vec_29[14];
    assign dep_chan_vld_29_16 = out_chan_dep_vld_vec_29[15];
    assign dep_chan_data_29_16 = out_chan_dep_data_29;
    assign token_29_16 = token_out_vec_29[15];
    assign dep_chan_vld_29_17 = out_chan_dep_vld_vec_29[16];
    assign dep_chan_data_29_17 = out_chan_dep_data_29;
    assign token_29_17 = token_out_vec_29[16];
    assign dep_chan_vld_29_18 = out_chan_dep_vld_vec_29[17];
    assign dep_chan_data_29_18 = out_chan_dep_data_29;
    assign token_29_18 = token_out_vec_29[17];
    assign dep_chan_vld_29_19 = out_chan_dep_vld_vec_29[18];
    assign dep_chan_data_29_19 = out_chan_dep_data_29;
    assign token_29_19 = token_out_vec_29[18];
    assign dep_chan_vld_29_20 = out_chan_dep_vld_vec_29[19];
    assign dep_chan_data_29_20 = out_chan_dep_data_29;
    assign token_29_20 = token_out_vec_29[19];
    assign dep_chan_vld_29_21 = out_chan_dep_vld_vec_29[20];
    assign dep_chan_data_29_21 = out_chan_dep_data_29;
    assign token_29_21 = token_out_vec_29[20];
    assign dep_chan_vld_29_22 = out_chan_dep_vld_vec_29[21];
    assign dep_chan_data_29_22 = out_chan_dep_data_29;
    assign token_29_22 = token_out_vec_29[21];
    assign dep_chan_vld_29_23 = out_chan_dep_vld_vec_29[22];
    assign dep_chan_data_29_23 = out_chan_dep_data_29;
    assign token_29_23 = token_out_vec_29[22];
    assign dep_chan_vld_29_24 = out_chan_dep_vld_vec_29[23];
    assign dep_chan_data_29_24 = out_chan_dep_data_29;
    assign token_29_24 = token_out_vec_29[23];
    assign dep_chan_vld_29_25 = out_chan_dep_vld_vec_29[24];
    assign dep_chan_data_29_25 = out_chan_dep_data_29;
    assign token_29_25 = token_out_vec_29[24];
    assign dep_chan_vld_29_26 = out_chan_dep_vld_vec_29[25];
    assign dep_chan_data_29_26 = out_chan_dep_data_29;
    assign token_29_26 = token_out_vec_29[25];
    assign dep_chan_vld_29_27 = out_chan_dep_vld_vec_29[26];
    assign dep_chan_data_29_27 = out_chan_dep_data_29;
    assign token_29_27 = token_out_vec_29[26];
    assign dep_chan_vld_29_31 = out_chan_dep_vld_vec_29[27];
    assign dep_chan_data_29_31 = out_chan_dep_data_29;
    assign token_29_31 = token_out_vec_29[27];
    assign dep_chan_vld_29_32 = out_chan_dep_vld_vec_29[28];
    assign dep_chan_data_29_32 = out_chan_dep_data_29;
    assign token_29_32 = token_out_vec_29[28];
    assign dep_chan_vld_29_33 = out_chan_dep_vld_vec_29[29];
    assign dep_chan_data_29_33 = out_chan_dep_data_29;
    assign token_29_33 = token_out_vec_29[29];
    assign dep_chan_vld_29_34 = out_chan_dep_vld_vec_29[30];
    assign dep_chan_data_29_34 = out_chan_dep_data_29;
    assign token_29_34 = token_out_vec_29[30];
    assign dep_chan_vld_29_35 = out_chan_dep_vld_vec_29[31];
    assign dep_chan_data_29_35 = out_chan_dep_data_29;
    assign token_29_35 = token_out_vec_29[31];
    assign dep_chan_vld_29_36 = out_chan_dep_vld_vec_29[32];
    assign dep_chan_data_29_36 = out_chan_dep_data_29;
    assign token_29_36 = token_out_vec_29[32];

    // Process: ProcessingElement_25_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 30, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_30 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_30),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_30),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_30),
        .token_in_vec(token_in_vec_30),
        .dl_detect_in(dl_detect_out),
        .origin(origin[30]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_30),
        .out_chan_dep_data(out_chan_dep_data_30),
        .token_out_vec(token_out_vec_30),
        .dl_detect_out(dl_in_vec[30]));

    assign proc_30_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_24_blk_n) | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_24_blk_n) | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_WriteC_Flattened_fu_179.cPipes_24_blk_n);
    assign proc_30_data_PIPO_blk[0] = 1'b0;
    assign proc_30_start_FIFO_blk[0] = 1'b0;
    assign proc_30_TLF_FIFO_blk[0] = 1'b0;
    assign proc_30_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_30_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_30[0] = dl_detect_out ? proc_dep_vld_vec_30_reg[0] : (proc_30_data_FIFO_blk[0] | proc_30_data_PIPO_blk[0] | proc_30_start_FIFO_blk[0] | proc_30_TLF_FIFO_blk[0] | proc_30_input_sync_blk[0] | proc_30_output_sync_blk[0]);
    assign proc_30_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_25_blk_n) | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_25_blk_n) | (~ProcessingElement_25_U0.grp_ProcessingElement_25_Pipeline_WriteC_Flattened_fu_179.cPipes_25_blk_n);
    assign proc_30_data_PIPO_blk[1] = 1'b0;
    assign proc_30_start_FIFO_blk[1] = 1'b0;
    assign proc_30_TLF_FIFO_blk[1] = 1'b0;
    assign proc_30_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_30_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_30[1] = dl_detect_out ? proc_dep_vld_vec_30_reg[1] : (proc_30_data_FIFO_blk[1] | proc_30_data_PIPO_blk[1] | proc_30_start_FIFO_blk[1] | proc_30_TLF_FIFO_blk[1] | proc_30_input_sync_blk[1] | proc_30_output_sync_blk[1]);
    assign proc_30_data_FIFO_blk[2] = 1'b0;
    assign proc_30_data_PIPO_blk[2] = 1'b0;
    assign proc_30_start_FIFO_blk[2] = 1'b0;
    assign proc_30_TLF_FIFO_blk[2] = 1'b0;
    assign proc_30_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_30_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_30[2] = dl_detect_out ? proc_dep_vld_vec_30_reg[2] : (proc_30_data_FIFO_blk[2] | proc_30_data_PIPO_blk[2] | proc_30_start_FIFO_blk[2] | proc_30_TLF_FIFO_blk[2] | proc_30_input_sync_blk[2] | proc_30_output_sync_blk[2]);
    assign proc_30_data_FIFO_blk[3] = 1'b0;
    assign proc_30_data_PIPO_blk[3] = 1'b0;
    assign proc_30_start_FIFO_blk[3] = 1'b0;
    assign proc_30_TLF_FIFO_blk[3] = 1'b0;
    assign proc_30_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_30_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_30[3] = dl_detect_out ? proc_dep_vld_vec_30_reg[3] : (proc_30_data_FIFO_blk[3] | proc_30_data_PIPO_blk[3] | proc_30_start_FIFO_blk[3] | proc_30_TLF_FIFO_blk[3] | proc_30_input_sync_blk[3] | proc_30_output_sync_blk[3]);
    assign proc_30_data_FIFO_blk[4] = 1'b0;
    assign proc_30_data_PIPO_blk[4] = 1'b0;
    assign proc_30_start_FIFO_blk[4] = 1'b0;
    assign proc_30_TLF_FIFO_blk[4] = 1'b0;
    assign proc_30_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_30_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_30[4] = dl_detect_out ? proc_dep_vld_vec_30_reg[4] : (proc_30_data_FIFO_blk[4] | proc_30_data_PIPO_blk[4] | proc_30_start_FIFO_blk[4] | proc_30_TLF_FIFO_blk[4] | proc_30_input_sync_blk[4] | proc_30_output_sync_blk[4]);
    assign proc_30_data_FIFO_blk[5] = 1'b0;
    assign proc_30_data_PIPO_blk[5] = 1'b0;
    assign proc_30_start_FIFO_blk[5] = 1'b0;
    assign proc_30_TLF_FIFO_blk[5] = 1'b0;
    assign proc_30_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_30_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_30[5] = dl_detect_out ? proc_dep_vld_vec_30_reg[5] : (proc_30_data_FIFO_blk[5] | proc_30_data_PIPO_blk[5] | proc_30_start_FIFO_blk[5] | proc_30_TLF_FIFO_blk[5] | proc_30_input_sync_blk[5] | proc_30_output_sync_blk[5]);
    assign proc_30_data_FIFO_blk[6] = 1'b0;
    assign proc_30_data_PIPO_blk[6] = 1'b0;
    assign proc_30_start_FIFO_blk[6] = 1'b0;
    assign proc_30_TLF_FIFO_blk[6] = 1'b0;
    assign proc_30_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_30_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_30[6] = dl_detect_out ? proc_dep_vld_vec_30_reg[6] : (proc_30_data_FIFO_blk[6] | proc_30_data_PIPO_blk[6] | proc_30_start_FIFO_blk[6] | proc_30_TLF_FIFO_blk[6] | proc_30_input_sync_blk[6] | proc_30_output_sync_blk[6]);
    assign proc_30_data_FIFO_blk[7] = 1'b0;
    assign proc_30_data_PIPO_blk[7] = 1'b0;
    assign proc_30_start_FIFO_blk[7] = 1'b0;
    assign proc_30_TLF_FIFO_blk[7] = 1'b0;
    assign proc_30_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_30_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_30[7] = dl_detect_out ? proc_dep_vld_vec_30_reg[7] : (proc_30_data_FIFO_blk[7] | proc_30_data_PIPO_blk[7] | proc_30_start_FIFO_blk[7] | proc_30_TLF_FIFO_blk[7] | proc_30_input_sync_blk[7] | proc_30_output_sync_blk[7]);
    assign proc_30_data_FIFO_blk[8] = 1'b0;
    assign proc_30_data_PIPO_blk[8] = 1'b0;
    assign proc_30_start_FIFO_blk[8] = 1'b0;
    assign proc_30_TLF_FIFO_blk[8] = 1'b0;
    assign proc_30_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_30_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_30[8] = dl_detect_out ? proc_dep_vld_vec_30_reg[8] : (proc_30_data_FIFO_blk[8] | proc_30_data_PIPO_blk[8] | proc_30_start_FIFO_blk[8] | proc_30_TLF_FIFO_blk[8] | proc_30_input_sync_blk[8] | proc_30_output_sync_blk[8]);
    assign proc_30_data_FIFO_blk[9] = 1'b0;
    assign proc_30_data_PIPO_blk[9] = 1'b0;
    assign proc_30_start_FIFO_blk[9] = 1'b0;
    assign proc_30_TLF_FIFO_blk[9] = 1'b0;
    assign proc_30_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_30_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_30[9] = dl_detect_out ? proc_dep_vld_vec_30_reg[9] : (proc_30_data_FIFO_blk[9] | proc_30_data_PIPO_blk[9] | proc_30_start_FIFO_blk[9] | proc_30_TLF_FIFO_blk[9] | proc_30_input_sync_blk[9] | proc_30_output_sync_blk[9]);
    assign proc_30_data_FIFO_blk[10] = 1'b0;
    assign proc_30_data_PIPO_blk[10] = 1'b0;
    assign proc_30_start_FIFO_blk[10] = 1'b0;
    assign proc_30_TLF_FIFO_blk[10] = 1'b0;
    assign proc_30_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_30_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_30[10] = dl_detect_out ? proc_dep_vld_vec_30_reg[10] : (proc_30_data_FIFO_blk[10] | proc_30_data_PIPO_blk[10] | proc_30_start_FIFO_blk[10] | proc_30_TLF_FIFO_blk[10] | proc_30_input_sync_blk[10] | proc_30_output_sync_blk[10]);
    assign proc_30_data_FIFO_blk[11] = 1'b0;
    assign proc_30_data_PIPO_blk[11] = 1'b0;
    assign proc_30_start_FIFO_blk[11] = 1'b0;
    assign proc_30_TLF_FIFO_blk[11] = 1'b0;
    assign proc_30_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_30_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_30[11] = dl_detect_out ? proc_dep_vld_vec_30_reg[11] : (proc_30_data_FIFO_blk[11] | proc_30_data_PIPO_blk[11] | proc_30_start_FIFO_blk[11] | proc_30_TLF_FIFO_blk[11] | proc_30_input_sync_blk[11] | proc_30_output_sync_blk[11]);
    assign proc_30_data_FIFO_blk[12] = 1'b0;
    assign proc_30_data_PIPO_blk[12] = 1'b0;
    assign proc_30_start_FIFO_blk[12] = 1'b0;
    assign proc_30_TLF_FIFO_blk[12] = 1'b0;
    assign proc_30_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_30_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_30[12] = dl_detect_out ? proc_dep_vld_vec_30_reg[12] : (proc_30_data_FIFO_blk[12] | proc_30_data_PIPO_blk[12] | proc_30_start_FIFO_blk[12] | proc_30_TLF_FIFO_blk[12] | proc_30_input_sync_blk[12] | proc_30_output_sync_blk[12]);
    assign proc_30_data_FIFO_blk[13] = 1'b0;
    assign proc_30_data_PIPO_blk[13] = 1'b0;
    assign proc_30_start_FIFO_blk[13] = 1'b0;
    assign proc_30_TLF_FIFO_blk[13] = 1'b0;
    assign proc_30_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_30_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_30[13] = dl_detect_out ? proc_dep_vld_vec_30_reg[13] : (proc_30_data_FIFO_blk[13] | proc_30_data_PIPO_blk[13] | proc_30_start_FIFO_blk[13] | proc_30_TLF_FIFO_blk[13] | proc_30_input_sync_blk[13] | proc_30_output_sync_blk[13]);
    assign proc_30_data_FIFO_blk[14] = 1'b0;
    assign proc_30_data_PIPO_blk[14] = 1'b0;
    assign proc_30_start_FIFO_blk[14] = 1'b0;
    assign proc_30_TLF_FIFO_blk[14] = 1'b0;
    assign proc_30_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_30_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_30[14] = dl_detect_out ? proc_dep_vld_vec_30_reg[14] : (proc_30_data_FIFO_blk[14] | proc_30_data_PIPO_blk[14] | proc_30_start_FIFO_blk[14] | proc_30_TLF_FIFO_blk[14] | proc_30_input_sync_blk[14] | proc_30_output_sync_blk[14]);
    assign proc_30_data_FIFO_blk[15] = 1'b0;
    assign proc_30_data_PIPO_blk[15] = 1'b0;
    assign proc_30_start_FIFO_blk[15] = 1'b0;
    assign proc_30_TLF_FIFO_blk[15] = 1'b0;
    assign proc_30_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_30_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_30[15] = dl_detect_out ? proc_dep_vld_vec_30_reg[15] : (proc_30_data_FIFO_blk[15] | proc_30_data_PIPO_blk[15] | proc_30_start_FIFO_blk[15] | proc_30_TLF_FIFO_blk[15] | proc_30_input_sync_blk[15] | proc_30_output_sync_blk[15]);
    assign proc_30_data_FIFO_blk[16] = 1'b0;
    assign proc_30_data_PIPO_blk[16] = 1'b0;
    assign proc_30_start_FIFO_blk[16] = 1'b0;
    assign proc_30_TLF_FIFO_blk[16] = 1'b0;
    assign proc_30_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_30_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_30[16] = dl_detect_out ? proc_dep_vld_vec_30_reg[16] : (proc_30_data_FIFO_blk[16] | proc_30_data_PIPO_blk[16] | proc_30_start_FIFO_blk[16] | proc_30_TLF_FIFO_blk[16] | proc_30_input_sync_blk[16] | proc_30_output_sync_blk[16]);
    assign proc_30_data_FIFO_blk[17] = 1'b0;
    assign proc_30_data_PIPO_blk[17] = 1'b0;
    assign proc_30_start_FIFO_blk[17] = 1'b0;
    assign proc_30_TLF_FIFO_blk[17] = 1'b0;
    assign proc_30_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_30_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_30[17] = dl_detect_out ? proc_dep_vld_vec_30_reg[17] : (proc_30_data_FIFO_blk[17] | proc_30_data_PIPO_blk[17] | proc_30_start_FIFO_blk[17] | proc_30_TLF_FIFO_blk[17] | proc_30_input_sync_blk[17] | proc_30_output_sync_blk[17]);
    assign proc_30_data_FIFO_blk[18] = 1'b0;
    assign proc_30_data_PIPO_blk[18] = 1'b0;
    assign proc_30_start_FIFO_blk[18] = 1'b0;
    assign proc_30_TLF_FIFO_blk[18] = 1'b0;
    assign proc_30_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_30_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_30[18] = dl_detect_out ? proc_dep_vld_vec_30_reg[18] : (proc_30_data_FIFO_blk[18] | proc_30_data_PIPO_blk[18] | proc_30_start_FIFO_blk[18] | proc_30_TLF_FIFO_blk[18] | proc_30_input_sync_blk[18] | proc_30_output_sync_blk[18]);
    assign proc_30_data_FIFO_blk[19] = 1'b0;
    assign proc_30_data_PIPO_blk[19] = 1'b0;
    assign proc_30_start_FIFO_blk[19] = 1'b0;
    assign proc_30_TLF_FIFO_blk[19] = 1'b0;
    assign proc_30_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_30_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_30[19] = dl_detect_out ? proc_dep_vld_vec_30_reg[19] : (proc_30_data_FIFO_blk[19] | proc_30_data_PIPO_blk[19] | proc_30_start_FIFO_blk[19] | proc_30_TLF_FIFO_blk[19] | proc_30_input_sync_blk[19] | proc_30_output_sync_blk[19]);
    assign proc_30_data_FIFO_blk[20] = 1'b0;
    assign proc_30_data_PIPO_blk[20] = 1'b0;
    assign proc_30_start_FIFO_blk[20] = 1'b0;
    assign proc_30_TLF_FIFO_blk[20] = 1'b0;
    assign proc_30_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_30_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_30[20] = dl_detect_out ? proc_dep_vld_vec_30_reg[20] : (proc_30_data_FIFO_blk[20] | proc_30_data_PIPO_blk[20] | proc_30_start_FIFO_blk[20] | proc_30_TLF_FIFO_blk[20] | proc_30_input_sync_blk[20] | proc_30_output_sync_blk[20]);
    assign proc_30_data_FIFO_blk[21] = 1'b0;
    assign proc_30_data_PIPO_blk[21] = 1'b0;
    assign proc_30_start_FIFO_blk[21] = 1'b0;
    assign proc_30_TLF_FIFO_blk[21] = 1'b0;
    assign proc_30_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_30_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_30[21] = dl_detect_out ? proc_dep_vld_vec_30_reg[21] : (proc_30_data_FIFO_blk[21] | proc_30_data_PIPO_blk[21] | proc_30_start_FIFO_blk[21] | proc_30_TLF_FIFO_blk[21] | proc_30_input_sync_blk[21] | proc_30_output_sync_blk[21]);
    assign proc_30_data_FIFO_blk[22] = 1'b0;
    assign proc_30_data_PIPO_blk[22] = 1'b0;
    assign proc_30_start_FIFO_blk[22] = 1'b0;
    assign proc_30_TLF_FIFO_blk[22] = 1'b0;
    assign proc_30_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_30_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_30[22] = dl_detect_out ? proc_dep_vld_vec_30_reg[22] : (proc_30_data_FIFO_blk[22] | proc_30_data_PIPO_blk[22] | proc_30_start_FIFO_blk[22] | proc_30_TLF_FIFO_blk[22] | proc_30_input_sync_blk[22] | proc_30_output_sync_blk[22]);
    assign proc_30_data_FIFO_blk[23] = 1'b0;
    assign proc_30_data_PIPO_blk[23] = 1'b0;
    assign proc_30_start_FIFO_blk[23] = 1'b0;
    assign proc_30_TLF_FIFO_blk[23] = 1'b0;
    assign proc_30_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_30_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_30[23] = dl_detect_out ? proc_dep_vld_vec_30_reg[23] : (proc_30_data_FIFO_blk[23] | proc_30_data_PIPO_blk[23] | proc_30_start_FIFO_blk[23] | proc_30_TLF_FIFO_blk[23] | proc_30_input_sync_blk[23] | proc_30_output_sync_blk[23]);
    assign proc_30_data_FIFO_blk[24] = 1'b0;
    assign proc_30_data_PIPO_blk[24] = 1'b0;
    assign proc_30_start_FIFO_blk[24] = 1'b0;
    assign proc_30_TLF_FIFO_blk[24] = 1'b0;
    assign proc_30_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_30_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_30[24] = dl_detect_out ? proc_dep_vld_vec_30_reg[24] : (proc_30_data_FIFO_blk[24] | proc_30_data_PIPO_blk[24] | proc_30_start_FIFO_blk[24] | proc_30_TLF_FIFO_blk[24] | proc_30_input_sync_blk[24] | proc_30_output_sync_blk[24]);
    assign proc_30_data_FIFO_blk[25] = 1'b0;
    assign proc_30_data_PIPO_blk[25] = 1'b0;
    assign proc_30_start_FIFO_blk[25] = 1'b0;
    assign proc_30_TLF_FIFO_blk[25] = 1'b0;
    assign proc_30_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_30_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_30[25] = dl_detect_out ? proc_dep_vld_vec_30_reg[25] : (proc_30_data_FIFO_blk[25] | proc_30_data_PIPO_blk[25] | proc_30_start_FIFO_blk[25] | proc_30_TLF_FIFO_blk[25] | proc_30_input_sync_blk[25] | proc_30_output_sync_blk[25]);
    assign proc_30_data_FIFO_blk[26] = 1'b0;
    assign proc_30_data_PIPO_blk[26] = 1'b0;
    assign proc_30_start_FIFO_blk[26] = 1'b0;
    assign proc_30_TLF_FIFO_blk[26] = 1'b0;
    assign proc_30_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_30_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_30[26] = dl_detect_out ? proc_dep_vld_vec_30_reg[26] : (proc_30_data_FIFO_blk[26] | proc_30_data_PIPO_blk[26] | proc_30_start_FIFO_blk[26] | proc_30_TLF_FIFO_blk[26] | proc_30_input_sync_blk[26] | proc_30_output_sync_blk[26]);
    assign proc_30_data_FIFO_blk[27] = 1'b0;
    assign proc_30_data_PIPO_blk[27] = 1'b0;
    assign proc_30_start_FIFO_blk[27] = 1'b0;
    assign proc_30_TLF_FIFO_blk[27] = 1'b0;
    assign proc_30_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_30_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_30[27] = dl_detect_out ? proc_dep_vld_vec_30_reg[27] : (proc_30_data_FIFO_blk[27] | proc_30_data_PIPO_blk[27] | proc_30_start_FIFO_blk[27] | proc_30_TLF_FIFO_blk[27] | proc_30_input_sync_blk[27] | proc_30_output_sync_blk[27]);
    assign proc_30_data_FIFO_blk[28] = 1'b0;
    assign proc_30_data_PIPO_blk[28] = 1'b0;
    assign proc_30_start_FIFO_blk[28] = 1'b0;
    assign proc_30_TLF_FIFO_blk[28] = 1'b0;
    assign proc_30_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_30_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_30[28] = dl_detect_out ? proc_dep_vld_vec_30_reg[28] : (proc_30_data_FIFO_blk[28] | proc_30_data_PIPO_blk[28] | proc_30_start_FIFO_blk[28] | proc_30_TLF_FIFO_blk[28] | proc_30_input_sync_blk[28] | proc_30_output_sync_blk[28]);
    assign proc_30_data_FIFO_blk[29] = 1'b0;
    assign proc_30_data_PIPO_blk[29] = 1'b0;
    assign proc_30_start_FIFO_blk[29] = 1'b0;
    assign proc_30_TLF_FIFO_blk[29] = 1'b0;
    assign proc_30_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_30_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_30[29] = dl_detect_out ? proc_dep_vld_vec_30_reg[29] : (proc_30_data_FIFO_blk[29] | proc_30_data_PIPO_blk[29] | proc_30_start_FIFO_blk[29] | proc_30_TLF_FIFO_blk[29] | proc_30_input_sync_blk[29] | proc_30_output_sync_blk[29]);
    assign proc_30_data_FIFO_blk[30] = 1'b0;
    assign proc_30_data_PIPO_blk[30] = 1'b0;
    assign proc_30_start_FIFO_blk[30] = 1'b0;
    assign proc_30_TLF_FIFO_blk[30] = 1'b0;
    assign proc_30_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_30_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_30[30] = dl_detect_out ? proc_dep_vld_vec_30_reg[30] : (proc_30_data_FIFO_blk[30] | proc_30_data_PIPO_blk[30] | proc_30_start_FIFO_blk[30] | proc_30_TLF_FIFO_blk[30] | proc_30_input_sync_blk[30] | proc_30_output_sync_blk[30]);
    assign proc_30_data_FIFO_blk[31] = 1'b0;
    assign proc_30_data_PIPO_blk[31] = 1'b0;
    assign proc_30_start_FIFO_blk[31] = 1'b0;
    assign proc_30_TLF_FIFO_blk[31] = 1'b0;
    assign proc_30_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_30_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_30[31] = dl_detect_out ? proc_dep_vld_vec_30_reg[31] : (proc_30_data_FIFO_blk[31] | proc_30_data_PIPO_blk[31] | proc_30_start_FIFO_blk[31] | proc_30_TLF_FIFO_blk[31] | proc_30_input_sync_blk[31] | proc_30_output_sync_blk[31]);
    assign proc_30_data_FIFO_blk[32] = 1'b0;
    assign proc_30_data_PIPO_blk[32] = 1'b0;
    assign proc_30_start_FIFO_blk[32] = 1'b0;
    assign proc_30_TLF_FIFO_blk[32] = 1'b0;
    assign proc_30_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_25_U0_ap_ready & ProcessingElement_25_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_30_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_30[32] = dl_detect_out ? proc_dep_vld_vec_30_reg[32] : (proc_30_data_FIFO_blk[32] | proc_30_data_PIPO_blk[32] | proc_30_start_FIFO_blk[32] | proc_30_TLF_FIFO_blk[32] | proc_30_input_sync_blk[32] | proc_30_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_30_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_30_reg <= proc_dep_vld_vec_30;
        end
    end
    assign in_chan_dep_vld_vec_30[0] = dep_chan_vld_0_30;
    assign in_chan_dep_data_vec_30[39 : 0] = dep_chan_data_0_30;
    assign token_in_vec_30[0] = token_0_30;
    assign in_chan_dep_vld_vec_30[1] = dep_chan_vld_1_30;
    assign in_chan_dep_data_vec_30[79 : 40] = dep_chan_data_1_30;
    assign token_in_vec_30[1] = token_1_30;
    assign in_chan_dep_vld_vec_30[2] = dep_chan_vld_3_30;
    assign in_chan_dep_data_vec_30[119 : 80] = dep_chan_data_3_30;
    assign token_in_vec_30[2] = token_3_30;
    assign in_chan_dep_vld_vec_30[3] = dep_chan_vld_6_30;
    assign in_chan_dep_data_vec_30[159 : 120] = dep_chan_data_6_30;
    assign token_in_vec_30[3] = token_6_30;
    assign in_chan_dep_vld_vec_30[4] = dep_chan_vld_7_30;
    assign in_chan_dep_data_vec_30[199 : 160] = dep_chan_data_7_30;
    assign token_in_vec_30[4] = token_7_30;
    assign in_chan_dep_vld_vec_30[5] = dep_chan_vld_8_30;
    assign in_chan_dep_data_vec_30[239 : 200] = dep_chan_data_8_30;
    assign token_in_vec_30[5] = token_8_30;
    assign in_chan_dep_vld_vec_30[6] = dep_chan_vld_9_30;
    assign in_chan_dep_data_vec_30[279 : 240] = dep_chan_data_9_30;
    assign token_in_vec_30[6] = token_9_30;
    assign in_chan_dep_vld_vec_30[7] = dep_chan_vld_10_30;
    assign in_chan_dep_data_vec_30[319 : 280] = dep_chan_data_10_30;
    assign token_in_vec_30[7] = token_10_30;
    assign in_chan_dep_vld_vec_30[8] = dep_chan_vld_11_30;
    assign in_chan_dep_data_vec_30[359 : 320] = dep_chan_data_11_30;
    assign token_in_vec_30[8] = token_11_30;
    assign in_chan_dep_vld_vec_30[9] = dep_chan_vld_12_30;
    assign in_chan_dep_data_vec_30[399 : 360] = dep_chan_data_12_30;
    assign token_in_vec_30[9] = token_12_30;
    assign in_chan_dep_vld_vec_30[10] = dep_chan_vld_13_30;
    assign in_chan_dep_data_vec_30[439 : 400] = dep_chan_data_13_30;
    assign token_in_vec_30[10] = token_13_30;
    assign in_chan_dep_vld_vec_30[11] = dep_chan_vld_14_30;
    assign in_chan_dep_data_vec_30[479 : 440] = dep_chan_data_14_30;
    assign token_in_vec_30[11] = token_14_30;
    assign in_chan_dep_vld_vec_30[12] = dep_chan_vld_15_30;
    assign in_chan_dep_data_vec_30[519 : 480] = dep_chan_data_15_30;
    assign token_in_vec_30[12] = token_15_30;
    assign in_chan_dep_vld_vec_30[13] = dep_chan_vld_16_30;
    assign in_chan_dep_data_vec_30[559 : 520] = dep_chan_data_16_30;
    assign token_in_vec_30[13] = token_16_30;
    assign in_chan_dep_vld_vec_30[14] = dep_chan_vld_17_30;
    assign in_chan_dep_data_vec_30[599 : 560] = dep_chan_data_17_30;
    assign token_in_vec_30[14] = token_17_30;
    assign in_chan_dep_vld_vec_30[15] = dep_chan_vld_18_30;
    assign in_chan_dep_data_vec_30[639 : 600] = dep_chan_data_18_30;
    assign token_in_vec_30[15] = token_18_30;
    assign in_chan_dep_vld_vec_30[16] = dep_chan_vld_19_30;
    assign in_chan_dep_data_vec_30[679 : 640] = dep_chan_data_19_30;
    assign token_in_vec_30[16] = token_19_30;
    assign in_chan_dep_vld_vec_30[17] = dep_chan_vld_20_30;
    assign in_chan_dep_data_vec_30[719 : 680] = dep_chan_data_20_30;
    assign token_in_vec_30[17] = token_20_30;
    assign in_chan_dep_vld_vec_30[18] = dep_chan_vld_21_30;
    assign in_chan_dep_data_vec_30[759 : 720] = dep_chan_data_21_30;
    assign token_in_vec_30[18] = token_21_30;
    assign in_chan_dep_vld_vec_30[19] = dep_chan_vld_22_30;
    assign in_chan_dep_data_vec_30[799 : 760] = dep_chan_data_22_30;
    assign token_in_vec_30[19] = token_22_30;
    assign in_chan_dep_vld_vec_30[20] = dep_chan_vld_23_30;
    assign in_chan_dep_data_vec_30[839 : 800] = dep_chan_data_23_30;
    assign token_in_vec_30[20] = token_23_30;
    assign in_chan_dep_vld_vec_30[21] = dep_chan_vld_24_30;
    assign in_chan_dep_data_vec_30[879 : 840] = dep_chan_data_24_30;
    assign token_in_vec_30[21] = token_24_30;
    assign in_chan_dep_vld_vec_30[22] = dep_chan_vld_25_30;
    assign in_chan_dep_data_vec_30[919 : 880] = dep_chan_data_25_30;
    assign token_in_vec_30[22] = token_25_30;
    assign in_chan_dep_vld_vec_30[23] = dep_chan_vld_26_30;
    assign in_chan_dep_data_vec_30[959 : 920] = dep_chan_data_26_30;
    assign token_in_vec_30[23] = token_26_30;
    assign in_chan_dep_vld_vec_30[24] = dep_chan_vld_27_30;
    assign in_chan_dep_data_vec_30[999 : 960] = dep_chan_data_27_30;
    assign token_in_vec_30[24] = token_27_30;
    assign in_chan_dep_vld_vec_30[25] = dep_chan_vld_28_30;
    assign in_chan_dep_data_vec_30[1039 : 1000] = dep_chan_data_28_30;
    assign token_in_vec_30[25] = token_28_30;
    assign in_chan_dep_vld_vec_30[26] = dep_chan_vld_29_30;
    assign in_chan_dep_data_vec_30[1079 : 1040] = dep_chan_data_29_30;
    assign token_in_vec_30[26] = token_29_30;
    assign in_chan_dep_vld_vec_30[27] = dep_chan_vld_31_30;
    assign in_chan_dep_data_vec_30[1119 : 1080] = dep_chan_data_31_30;
    assign token_in_vec_30[27] = token_31_30;
    assign in_chan_dep_vld_vec_30[28] = dep_chan_vld_32_30;
    assign in_chan_dep_data_vec_30[1159 : 1120] = dep_chan_data_32_30;
    assign token_in_vec_30[28] = token_32_30;
    assign in_chan_dep_vld_vec_30[29] = dep_chan_vld_33_30;
    assign in_chan_dep_data_vec_30[1199 : 1160] = dep_chan_data_33_30;
    assign token_in_vec_30[29] = token_33_30;
    assign in_chan_dep_vld_vec_30[30] = dep_chan_vld_34_30;
    assign in_chan_dep_data_vec_30[1239 : 1200] = dep_chan_data_34_30;
    assign token_in_vec_30[30] = token_34_30;
    assign in_chan_dep_vld_vec_30[31] = dep_chan_vld_35_30;
    assign in_chan_dep_data_vec_30[1279 : 1240] = dep_chan_data_35_30;
    assign token_in_vec_30[31] = token_35_30;
    assign in_chan_dep_vld_vec_30[32] = dep_chan_vld_36_30;
    assign in_chan_dep_data_vec_30[1319 : 1280] = dep_chan_data_36_30;
    assign token_in_vec_30[32] = token_36_30;
    assign dep_chan_vld_30_29 = out_chan_dep_vld_vec_30[0];
    assign dep_chan_data_30_29 = out_chan_dep_data_30;
    assign token_30_29 = token_out_vec_30[0];
    assign dep_chan_vld_30_31 = out_chan_dep_vld_vec_30[1];
    assign dep_chan_data_30_31 = out_chan_dep_data_30;
    assign token_30_31 = token_out_vec_30[1];
    assign dep_chan_vld_30_0 = out_chan_dep_vld_vec_30[2];
    assign dep_chan_data_30_0 = out_chan_dep_data_30;
    assign token_30_0 = token_out_vec_30[2];
    assign dep_chan_vld_30_1 = out_chan_dep_vld_vec_30[3];
    assign dep_chan_data_30_1 = out_chan_dep_data_30;
    assign token_30_1 = token_out_vec_30[3];
    assign dep_chan_vld_30_3 = out_chan_dep_vld_vec_30[4];
    assign dep_chan_data_30_3 = out_chan_dep_data_30;
    assign token_30_3 = token_out_vec_30[4];
    assign dep_chan_vld_30_6 = out_chan_dep_vld_vec_30[5];
    assign dep_chan_data_30_6 = out_chan_dep_data_30;
    assign token_30_6 = token_out_vec_30[5];
    assign dep_chan_vld_30_7 = out_chan_dep_vld_vec_30[6];
    assign dep_chan_data_30_7 = out_chan_dep_data_30;
    assign token_30_7 = token_out_vec_30[6];
    assign dep_chan_vld_30_8 = out_chan_dep_vld_vec_30[7];
    assign dep_chan_data_30_8 = out_chan_dep_data_30;
    assign token_30_8 = token_out_vec_30[7];
    assign dep_chan_vld_30_9 = out_chan_dep_vld_vec_30[8];
    assign dep_chan_data_30_9 = out_chan_dep_data_30;
    assign token_30_9 = token_out_vec_30[8];
    assign dep_chan_vld_30_10 = out_chan_dep_vld_vec_30[9];
    assign dep_chan_data_30_10 = out_chan_dep_data_30;
    assign token_30_10 = token_out_vec_30[9];
    assign dep_chan_vld_30_11 = out_chan_dep_vld_vec_30[10];
    assign dep_chan_data_30_11 = out_chan_dep_data_30;
    assign token_30_11 = token_out_vec_30[10];
    assign dep_chan_vld_30_12 = out_chan_dep_vld_vec_30[11];
    assign dep_chan_data_30_12 = out_chan_dep_data_30;
    assign token_30_12 = token_out_vec_30[11];
    assign dep_chan_vld_30_13 = out_chan_dep_vld_vec_30[12];
    assign dep_chan_data_30_13 = out_chan_dep_data_30;
    assign token_30_13 = token_out_vec_30[12];
    assign dep_chan_vld_30_14 = out_chan_dep_vld_vec_30[13];
    assign dep_chan_data_30_14 = out_chan_dep_data_30;
    assign token_30_14 = token_out_vec_30[13];
    assign dep_chan_vld_30_15 = out_chan_dep_vld_vec_30[14];
    assign dep_chan_data_30_15 = out_chan_dep_data_30;
    assign token_30_15 = token_out_vec_30[14];
    assign dep_chan_vld_30_16 = out_chan_dep_vld_vec_30[15];
    assign dep_chan_data_30_16 = out_chan_dep_data_30;
    assign token_30_16 = token_out_vec_30[15];
    assign dep_chan_vld_30_17 = out_chan_dep_vld_vec_30[16];
    assign dep_chan_data_30_17 = out_chan_dep_data_30;
    assign token_30_17 = token_out_vec_30[16];
    assign dep_chan_vld_30_18 = out_chan_dep_vld_vec_30[17];
    assign dep_chan_data_30_18 = out_chan_dep_data_30;
    assign token_30_18 = token_out_vec_30[17];
    assign dep_chan_vld_30_19 = out_chan_dep_vld_vec_30[18];
    assign dep_chan_data_30_19 = out_chan_dep_data_30;
    assign token_30_19 = token_out_vec_30[18];
    assign dep_chan_vld_30_20 = out_chan_dep_vld_vec_30[19];
    assign dep_chan_data_30_20 = out_chan_dep_data_30;
    assign token_30_20 = token_out_vec_30[19];
    assign dep_chan_vld_30_21 = out_chan_dep_vld_vec_30[20];
    assign dep_chan_data_30_21 = out_chan_dep_data_30;
    assign token_30_21 = token_out_vec_30[20];
    assign dep_chan_vld_30_22 = out_chan_dep_vld_vec_30[21];
    assign dep_chan_data_30_22 = out_chan_dep_data_30;
    assign token_30_22 = token_out_vec_30[21];
    assign dep_chan_vld_30_23 = out_chan_dep_vld_vec_30[22];
    assign dep_chan_data_30_23 = out_chan_dep_data_30;
    assign token_30_23 = token_out_vec_30[22];
    assign dep_chan_vld_30_24 = out_chan_dep_vld_vec_30[23];
    assign dep_chan_data_30_24 = out_chan_dep_data_30;
    assign token_30_24 = token_out_vec_30[23];
    assign dep_chan_vld_30_25 = out_chan_dep_vld_vec_30[24];
    assign dep_chan_data_30_25 = out_chan_dep_data_30;
    assign token_30_25 = token_out_vec_30[24];
    assign dep_chan_vld_30_26 = out_chan_dep_vld_vec_30[25];
    assign dep_chan_data_30_26 = out_chan_dep_data_30;
    assign token_30_26 = token_out_vec_30[25];
    assign dep_chan_vld_30_27 = out_chan_dep_vld_vec_30[26];
    assign dep_chan_data_30_27 = out_chan_dep_data_30;
    assign token_30_27 = token_out_vec_30[26];
    assign dep_chan_vld_30_28 = out_chan_dep_vld_vec_30[27];
    assign dep_chan_data_30_28 = out_chan_dep_data_30;
    assign token_30_28 = token_out_vec_30[27];
    assign dep_chan_vld_30_32 = out_chan_dep_vld_vec_30[28];
    assign dep_chan_data_30_32 = out_chan_dep_data_30;
    assign token_30_32 = token_out_vec_30[28];
    assign dep_chan_vld_30_33 = out_chan_dep_vld_vec_30[29];
    assign dep_chan_data_30_33 = out_chan_dep_data_30;
    assign token_30_33 = token_out_vec_30[29];
    assign dep_chan_vld_30_34 = out_chan_dep_vld_vec_30[30];
    assign dep_chan_data_30_34 = out_chan_dep_data_30;
    assign token_30_34 = token_out_vec_30[30];
    assign dep_chan_vld_30_35 = out_chan_dep_vld_vec_30[31];
    assign dep_chan_data_30_35 = out_chan_dep_data_30;
    assign token_30_35 = token_out_vec_30[31];
    assign dep_chan_vld_30_36 = out_chan_dep_vld_vec_30[32];
    assign dep_chan_data_30_36 = out_chan_dep_data_30;
    assign token_30_36 = token_out_vec_30[32];

    // Process: ProcessingElement_26_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 31, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_31 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_31),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_31),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_31),
        .token_in_vec(token_in_vec_31),
        .dl_detect_in(dl_detect_out),
        .origin(origin[31]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_31),
        .out_chan_dep_data(out_chan_dep_data_31),
        .token_out_vec(token_out_vec_31),
        .dl_detect_out(dl_in_vec[31]));

    assign proc_31_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_25_blk_n) | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_25_blk_n) | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_WriteC_Flattened_fu_179.cPipes_25_blk_n);
    assign proc_31_data_PIPO_blk[0] = 1'b0;
    assign proc_31_start_FIFO_blk[0] = 1'b0;
    assign proc_31_TLF_FIFO_blk[0] = 1'b0;
    assign proc_31_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_31_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_31[0] = dl_detect_out ? proc_dep_vld_vec_31_reg[0] : (proc_31_data_FIFO_blk[0] | proc_31_data_PIPO_blk[0] | proc_31_start_FIFO_blk[0] | proc_31_TLF_FIFO_blk[0] | proc_31_input_sync_blk[0] | proc_31_output_sync_blk[0]);
    assign proc_31_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_26_blk_n) | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_26_blk_n) | (~ProcessingElement_26_U0.grp_ProcessingElement_26_Pipeline_WriteC_Flattened_fu_179.cPipes_26_blk_n);
    assign proc_31_data_PIPO_blk[1] = 1'b0;
    assign proc_31_start_FIFO_blk[1] = 1'b0;
    assign proc_31_TLF_FIFO_blk[1] = 1'b0;
    assign proc_31_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_31_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_31[1] = dl_detect_out ? proc_dep_vld_vec_31_reg[1] : (proc_31_data_FIFO_blk[1] | proc_31_data_PIPO_blk[1] | proc_31_start_FIFO_blk[1] | proc_31_TLF_FIFO_blk[1] | proc_31_input_sync_blk[1] | proc_31_output_sync_blk[1]);
    assign proc_31_data_FIFO_blk[2] = 1'b0;
    assign proc_31_data_PIPO_blk[2] = 1'b0;
    assign proc_31_start_FIFO_blk[2] = 1'b0;
    assign proc_31_TLF_FIFO_blk[2] = 1'b0;
    assign proc_31_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_31_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_31[2] = dl_detect_out ? proc_dep_vld_vec_31_reg[2] : (proc_31_data_FIFO_blk[2] | proc_31_data_PIPO_blk[2] | proc_31_start_FIFO_blk[2] | proc_31_TLF_FIFO_blk[2] | proc_31_input_sync_blk[2] | proc_31_output_sync_blk[2]);
    assign proc_31_data_FIFO_blk[3] = 1'b0;
    assign proc_31_data_PIPO_blk[3] = 1'b0;
    assign proc_31_start_FIFO_blk[3] = 1'b0;
    assign proc_31_TLF_FIFO_blk[3] = 1'b0;
    assign proc_31_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_31_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_31[3] = dl_detect_out ? proc_dep_vld_vec_31_reg[3] : (proc_31_data_FIFO_blk[3] | proc_31_data_PIPO_blk[3] | proc_31_start_FIFO_blk[3] | proc_31_TLF_FIFO_blk[3] | proc_31_input_sync_blk[3] | proc_31_output_sync_blk[3]);
    assign proc_31_data_FIFO_blk[4] = 1'b0;
    assign proc_31_data_PIPO_blk[4] = 1'b0;
    assign proc_31_start_FIFO_blk[4] = 1'b0;
    assign proc_31_TLF_FIFO_blk[4] = 1'b0;
    assign proc_31_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_31_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_31[4] = dl_detect_out ? proc_dep_vld_vec_31_reg[4] : (proc_31_data_FIFO_blk[4] | proc_31_data_PIPO_blk[4] | proc_31_start_FIFO_blk[4] | proc_31_TLF_FIFO_blk[4] | proc_31_input_sync_blk[4] | proc_31_output_sync_blk[4]);
    assign proc_31_data_FIFO_blk[5] = 1'b0;
    assign proc_31_data_PIPO_blk[5] = 1'b0;
    assign proc_31_start_FIFO_blk[5] = 1'b0;
    assign proc_31_TLF_FIFO_blk[5] = 1'b0;
    assign proc_31_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_31_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_31[5] = dl_detect_out ? proc_dep_vld_vec_31_reg[5] : (proc_31_data_FIFO_blk[5] | proc_31_data_PIPO_blk[5] | proc_31_start_FIFO_blk[5] | proc_31_TLF_FIFO_blk[5] | proc_31_input_sync_blk[5] | proc_31_output_sync_blk[5]);
    assign proc_31_data_FIFO_blk[6] = 1'b0;
    assign proc_31_data_PIPO_blk[6] = 1'b0;
    assign proc_31_start_FIFO_blk[6] = 1'b0;
    assign proc_31_TLF_FIFO_blk[6] = 1'b0;
    assign proc_31_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_31_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_31[6] = dl_detect_out ? proc_dep_vld_vec_31_reg[6] : (proc_31_data_FIFO_blk[6] | proc_31_data_PIPO_blk[6] | proc_31_start_FIFO_blk[6] | proc_31_TLF_FIFO_blk[6] | proc_31_input_sync_blk[6] | proc_31_output_sync_blk[6]);
    assign proc_31_data_FIFO_blk[7] = 1'b0;
    assign proc_31_data_PIPO_blk[7] = 1'b0;
    assign proc_31_start_FIFO_blk[7] = 1'b0;
    assign proc_31_TLF_FIFO_blk[7] = 1'b0;
    assign proc_31_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_31_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_31[7] = dl_detect_out ? proc_dep_vld_vec_31_reg[7] : (proc_31_data_FIFO_blk[7] | proc_31_data_PIPO_blk[7] | proc_31_start_FIFO_blk[7] | proc_31_TLF_FIFO_blk[7] | proc_31_input_sync_blk[7] | proc_31_output_sync_blk[7]);
    assign proc_31_data_FIFO_blk[8] = 1'b0;
    assign proc_31_data_PIPO_blk[8] = 1'b0;
    assign proc_31_start_FIFO_blk[8] = 1'b0;
    assign proc_31_TLF_FIFO_blk[8] = 1'b0;
    assign proc_31_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_31_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_31[8] = dl_detect_out ? proc_dep_vld_vec_31_reg[8] : (proc_31_data_FIFO_blk[8] | proc_31_data_PIPO_blk[8] | proc_31_start_FIFO_blk[8] | proc_31_TLF_FIFO_blk[8] | proc_31_input_sync_blk[8] | proc_31_output_sync_blk[8]);
    assign proc_31_data_FIFO_blk[9] = 1'b0;
    assign proc_31_data_PIPO_blk[9] = 1'b0;
    assign proc_31_start_FIFO_blk[9] = 1'b0;
    assign proc_31_TLF_FIFO_blk[9] = 1'b0;
    assign proc_31_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_31_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_31[9] = dl_detect_out ? proc_dep_vld_vec_31_reg[9] : (proc_31_data_FIFO_blk[9] | proc_31_data_PIPO_blk[9] | proc_31_start_FIFO_blk[9] | proc_31_TLF_FIFO_blk[9] | proc_31_input_sync_blk[9] | proc_31_output_sync_blk[9]);
    assign proc_31_data_FIFO_blk[10] = 1'b0;
    assign proc_31_data_PIPO_blk[10] = 1'b0;
    assign proc_31_start_FIFO_blk[10] = 1'b0;
    assign proc_31_TLF_FIFO_blk[10] = 1'b0;
    assign proc_31_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_31_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_31[10] = dl_detect_out ? proc_dep_vld_vec_31_reg[10] : (proc_31_data_FIFO_blk[10] | proc_31_data_PIPO_blk[10] | proc_31_start_FIFO_blk[10] | proc_31_TLF_FIFO_blk[10] | proc_31_input_sync_blk[10] | proc_31_output_sync_blk[10]);
    assign proc_31_data_FIFO_blk[11] = 1'b0;
    assign proc_31_data_PIPO_blk[11] = 1'b0;
    assign proc_31_start_FIFO_blk[11] = 1'b0;
    assign proc_31_TLF_FIFO_blk[11] = 1'b0;
    assign proc_31_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_31_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_31[11] = dl_detect_out ? proc_dep_vld_vec_31_reg[11] : (proc_31_data_FIFO_blk[11] | proc_31_data_PIPO_blk[11] | proc_31_start_FIFO_blk[11] | proc_31_TLF_FIFO_blk[11] | proc_31_input_sync_blk[11] | proc_31_output_sync_blk[11]);
    assign proc_31_data_FIFO_blk[12] = 1'b0;
    assign proc_31_data_PIPO_blk[12] = 1'b0;
    assign proc_31_start_FIFO_blk[12] = 1'b0;
    assign proc_31_TLF_FIFO_blk[12] = 1'b0;
    assign proc_31_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_31_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_31[12] = dl_detect_out ? proc_dep_vld_vec_31_reg[12] : (proc_31_data_FIFO_blk[12] | proc_31_data_PIPO_blk[12] | proc_31_start_FIFO_blk[12] | proc_31_TLF_FIFO_blk[12] | proc_31_input_sync_blk[12] | proc_31_output_sync_blk[12]);
    assign proc_31_data_FIFO_blk[13] = 1'b0;
    assign proc_31_data_PIPO_blk[13] = 1'b0;
    assign proc_31_start_FIFO_blk[13] = 1'b0;
    assign proc_31_TLF_FIFO_blk[13] = 1'b0;
    assign proc_31_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_31_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_31[13] = dl_detect_out ? proc_dep_vld_vec_31_reg[13] : (proc_31_data_FIFO_blk[13] | proc_31_data_PIPO_blk[13] | proc_31_start_FIFO_blk[13] | proc_31_TLF_FIFO_blk[13] | proc_31_input_sync_blk[13] | proc_31_output_sync_blk[13]);
    assign proc_31_data_FIFO_blk[14] = 1'b0;
    assign proc_31_data_PIPO_blk[14] = 1'b0;
    assign proc_31_start_FIFO_blk[14] = 1'b0;
    assign proc_31_TLF_FIFO_blk[14] = 1'b0;
    assign proc_31_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_31_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_31[14] = dl_detect_out ? proc_dep_vld_vec_31_reg[14] : (proc_31_data_FIFO_blk[14] | proc_31_data_PIPO_blk[14] | proc_31_start_FIFO_blk[14] | proc_31_TLF_FIFO_blk[14] | proc_31_input_sync_blk[14] | proc_31_output_sync_blk[14]);
    assign proc_31_data_FIFO_blk[15] = 1'b0;
    assign proc_31_data_PIPO_blk[15] = 1'b0;
    assign proc_31_start_FIFO_blk[15] = 1'b0;
    assign proc_31_TLF_FIFO_blk[15] = 1'b0;
    assign proc_31_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_31_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_31[15] = dl_detect_out ? proc_dep_vld_vec_31_reg[15] : (proc_31_data_FIFO_blk[15] | proc_31_data_PIPO_blk[15] | proc_31_start_FIFO_blk[15] | proc_31_TLF_FIFO_blk[15] | proc_31_input_sync_blk[15] | proc_31_output_sync_blk[15]);
    assign proc_31_data_FIFO_blk[16] = 1'b0;
    assign proc_31_data_PIPO_blk[16] = 1'b0;
    assign proc_31_start_FIFO_blk[16] = 1'b0;
    assign proc_31_TLF_FIFO_blk[16] = 1'b0;
    assign proc_31_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_31_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_31[16] = dl_detect_out ? proc_dep_vld_vec_31_reg[16] : (proc_31_data_FIFO_blk[16] | proc_31_data_PIPO_blk[16] | proc_31_start_FIFO_blk[16] | proc_31_TLF_FIFO_blk[16] | proc_31_input_sync_blk[16] | proc_31_output_sync_blk[16]);
    assign proc_31_data_FIFO_blk[17] = 1'b0;
    assign proc_31_data_PIPO_blk[17] = 1'b0;
    assign proc_31_start_FIFO_blk[17] = 1'b0;
    assign proc_31_TLF_FIFO_blk[17] = 1'b0;
    assign proc_31_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_31_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_31[17] = dl_detect_out ? proc_dep_vld_vec_31_reg[17] : (proc_31_data_FIFO_blk[17] | proc_31_data_PIPO_blk[17] | proc_31_start_FIFO_blk[17] | proc_31_TLF_FIFO_blk[17] | proc_31_input_sync_blk[17] | proc_31_output_sync_blk[17]);
    assign proc_31_data_FIFO_blk[18] = 1'b0;
    assign proc_31_data_PIPO_blk[18] = 1'b0;
    assign proc_31_start_FIFO_blk[18] = 1'b0;
    assign proc_31_TLF_FIFO_blk[18] = 1'b0;
    assign proc_31_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_31_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_31[18] = dl_detect_out ? proc_dep_vld_vec_31_reg[18] : (proc_31_data_FIFO_blk[18] | proc_31_data_PIPO_blk[18] | proc_31_start_FIFO_blk[18] | proc_31_TLF_FIFO_blk[18] | proc_31_input_sync_blk[18] | proc_31_output_sync_blk[18]);
    assign proc_31_data_FIFO_blk[19] = 1'b0;
    assign proc_31_data_PIPO_blk[19] = 1'b0;
    assign proc_31_start_FIFO_blk[19] = 1'b0;
    assign proc_31_TLF_FIFO_blk[19] = 1'b0;
    assign proc_31_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_31_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_31[19] = dl_detect_out ? proc_dep_vld_vec_31_reg[19] : (proc_31_data_FIFO_blk[19] | proc_31_data_PIPO_blk[19] | proc_31_start_FIFO_blk[19] | proc_31_TLF_FIFO_blk[19] | proc_31_input_sync_blk[19] | proc_31_output_sync_blk[19]);
    assign proc_31_data_FIFO_blk[20] = 1'b0;
    assign proc_31_data_PIPO_blk[20] = 1'b0;
    assign proc_31_start_FIFO_blk[20] = 1'b0;
    assign proc_31_TLF_FIFO_blk[20] = 1'b0;
    assign proc_31_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_31_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_31[20] = dl_detect_out ? proc_dep_vld_vec_31_reg[20] : (proc_31_data_FIFO_blk[20] | proc_31_data_PIPO_blk[20] | proc_31_start_FIFO_blk[20] | proc_31_TLF_FIFO_blk[20] | proc_31_input_sync_blk[20] | proc_31_output_sync_blk[20]);
    assign proc_31_data_FIFO_blk[21] = 1'b0;
    assign proc_31_data_PIPO_blk[21] = 1'b0;
    assign proc_31_start_FIFO_blk[21] = 1'b0;
    assign proc_31_TLF_FIFO_blk[21] = 1'b0;
    assign proc_31_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_31_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_31[21] = dl_detect_out ? proc_dep_vld_vec_31_reg[21] : (proc_31_data_FIFO_blk[21] | proc_31_data_PIPO_blk[21] | proc_31_start_FIFO_blk[21] | proc_31_TLF_FIFO_blk[21] | proc_31_input_sync_blk[21] | proc_31_output_sync_blk[21]);
    assign proc_31_data_FIFO_blk[22] = 1'b0;
    assign proc_31_data_PIPO_blk[22] = 1'b0;
    assign proc_31_start_FIFO_blk[22] = 1'b0;
    assign proc_31_TLF_FIFO_blk[22] = 1'b0;
    assign proc_31_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_31_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_31[22] = dl_detect_out ? proc_dep_vld_vec_31_reg[22] : (proc_31_data_FIFO_blk[22] | proc_31_data_PIPO_blk[22] | proc_31_start_FIFO_blk[22] | proc_31_TLF_FIFO_blk[22] | proc_31_input_sync_blk[22] | proc_31_output_sync_blk[22]);
    assign proc_31_data_FIFO_blk[23] = 1'b0;
    assign proc_31_data_PIPO_blk[23] = 1'b0;
    assign proc_31_start_FIFO_blk[23] = 1'b0;
    assign proc_31_TLF_FIFO_blk[23] = 1'b0;
    assign proc_31_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_31_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_31[23] = dl_detect_out ? proc_dep_vld_vec_31_reg[23] : (proc_31_data_FIFO_blk[23] | proc_31_data_PIPO_blk[23] | proc_31_start_FIFO_blk[23] | proc_31_TLF_FIFO_blk[23] | proc_31_input_sync_blk[23] | proc_31_output_sync_blk[23]);
    assign proc_31_data_FIFO_blk[24] = 1'b0;
    assign proc_31_data_PIPO_blk[24] = 1'b0;
    assign proc_31_start_FIFO_blk[24] = 1'b0;
    assign proc_31_TLF_FIFO_blk[24] = 1'b0;
    assign proc_31_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_31_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_31[24] = dl_detect_out ? proc_dep_vld_vec_31_reg[24] : (proc_31_data_FIFO_blk[24] | proc_31_data_PIPO_blk[24] | proc_31_start_FIFO_blk[24] | proc_31_TLF_FIFO_blk[24] | proc_31_input_sync_blk[24] | proc_31_output_sync_blk[24]);
    assign proc_31_data_FIFO_blk[25] = 1'b0;
    assign proc_31_data_PIPO_blk[25] = 1'b0;
    assign proc_31_start_FIFO_blk[25] = 1'b0;
    assign proc_31_TLF_FIFO_blk[25] = 1'b0;
    assign proc_31_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_31_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_31[25] = dl_detect_out ? proc_dep_vld_vec_31_reg[25] : (proc_31_data_FIFO_blk[25] | proc_31_data_PIPO_blk[25] | proc_31_start_FIFO_blk[25] | proc_31_TLF_FIFO_blk[25] | proc_31_input_sync_blk[25] | proc_31_output_sync_blk[25]);
    assign proc_31_data_FIFO_blk[26] = 1'b0;
    assign proc_31_data_PIPO_blk[26] = 1'b0;
    assign proc_31_start_FIFO_blk[26] = 1'b0;
    assign proc_31_TLF_FIFO_blk[26] = 1'b0;
    assign proc_31_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_31_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_31[26] = dl_detect_out ? proc_dep_vld_vec_31_reg[26] : (proc_31_data_FIFO_blk[26] | proc_31_data_PIPO_blk[26] | proc_31_start_FIFO_blk[26] | proc_31_TLF_FIFO_blk[26] | proc_31_input_sync_blk[26] | proc_31_output_sync_blk[26]);
    assign proc_31_data_FIFO_blk[27] = 1'b0;
    assign proc_31_data_PIPO_blk[27] = 1'b0;
    assign proc_31_start_FIFO_blk[27] = 1'b0;
    assign proc_31_TLF_FIFO_blk[27] = 1'b0;
    assign proc_31_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_31_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_31[27] = dl_detect_out ? proc_dep_vld_vec_31_reg[27] : (proc_31_data_FIFO_blk[27] | proc_31_data_PIPO_blk[27] | proc_31_start_FIFO_blk[27] | proc_31_TLF_FIFO_blk[27] | proc_31_input_sync_blk[27] | proc_31_output_sync_blk[27]);
    assign proc_31_data_FIFO_blk[28] = 1'b0;
    assign proc_31_data_PIPO_blk[28] = 1'b0;
    assign proc_31_start_FIFO_blk[28] = 1'b0;
    assign proc_31_TLF_FIFO_blk[28] = 1'b0;
    assign proc_31_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_31_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_31[28] = dl_detect_out ? proc_dep_vld_vec_31_reg[28] : (proc_31_data_FIFO_blk[28] | proc_31_data_PIPO_blk[28] | proc_31_start_FIFO_blk[28] | proc_31_TLF_FIFO_blk[28] | proc_31_input_sync_blk[28] | proc_31_output_sync_blk[28]);
    assign proc_31_data_FIFO_blk[29] = 1'b0;
    assign proc_31_data_PIPO_blk[29] = 1'b0;
    assign proc_31_start_FIFO_blk[29] = 1'b0;
    assign proc_31_TLF_FIFO_blk[29] = 1'b0;
    assign proc_31_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_31_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_31[29] = dl_detect_out ? proc_dep_vld_vec_31_reg[29] : (proc_31_data_FIFO_blk[29] | proc_31_data_PIPO_blk[29] | proc_31_start_FIFO_blk[29] | proc_31_TLF_FIFO_blk[29] | proc_31_input_sync_blk[29] | proc_31_output_sync_blk[29]);
    assign proc_31_data_FIFO_blk[30] = 1'b0;
    assign proc_31_data_PIPO_blk[30] = 1'b0;
    assign proc_31_start_FIFO_blk[30] = 1'b0;
    assign proc_31_TLF_FIFO_blk[30] = 1'b0;
    assign proc_31_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_31_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_31[30] = dl_detect_out ? proc_dep_vld_vec_31_reg[30] : (proc_31_data_FIFO_blk[30] | proc_31_data_PIPO_blk[30] | proc_31_start_FIFO_blk[30] | proc_31_TLF_FIFO_blk[30] | proc_31_input_sync_blk[30] | proc_31_output_sync_blk[30]);
    assign proc_31_data_FIFO_blk[31] = 1'b0;
    assign proc_31_data_PIPO_blk[31] = 1'b0;
    assign proc_31_start_FIFO_blk[31] = 1'b0;
    assign proc_31_TLF_FIFO_blk[31] = 1'b0;
    assign proc_31_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_31_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_31[31] = dl_detect_out ? proc_dep_vld_vec_31_reg[31] : (proc_31_data_FIFO_blk[31] | proc_31_data_PIPO_blk[31] | proc_31_start_FIFO_blk[31] | proc_31_TLF_FIFO_blk[31] | proc_31_input_sync_blk[31] | proc_31_output_sync_blk[31]);
    assign proc_31_data_FIFO_blk[32] = 1'b0;
    assign proc_31_data_PIPO_blk[32] = 1'b0;
    assign proc_31_start_FIFO_blk[32] = 1'b0;
    assign proc_31_TLF_FIFO_blk[32] = 1'b0;
    assign proc_31_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_26_U0_ap_ready & ProcessingElement_26_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_31_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_31[32] = dl_detect_out ? proc_dep_vld_vec_31_reg[32] : (proc_31_data_FIFO_blk[32] | proc_31_data_PIPO_blk[32] | proc_31_start_FIFO_blk[32] | proc_31_TLF_FIFO_blk[32] | proc_31_input_sync_blk[32] | proc_31_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_31_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_31_reg <= proc_dep_vld_vec_31;
        end
    end
    assign in_chan_dep_vld_vec_31[0] = dep_chan_vld_0_31;
    assign in_chan_dep_data_vec_31[39 : 0] = dep_chan_data_0_31;
    assign token_in_vec_31[0] = token_0_31;
    assign in_chan_dep_vld_vec_31[1] = dep_chan_vld_1_31;
    assign in_chan_dep_data_vec_31[79 : 40] = dep_chan_data_1_31;
    assign token_in_vec_31[1] = token_1_31;
    assign in_chan_dep_vld_vec_31[2] = dep_chan_vld_3_31;
    assign in_chan_dep_data_vec_31[119 : 80] = dep_chan_data_3_31;
    assign token_in_vec_31[2] = token_3_31;
    assign in_chan_dep_vld_vec_31[3] = dep_chan_vld_6_31;
    assign in_chan_dep_data_vec_31[159 : 120] = dep_chan_data_6_31;
    assign token_in_vec_31[3] = token_6_31;
    assign in_chan_dep_vld_vec_31[4] = dep_chan_vld_7_31;
    assign in_chan_dep_data_vec_31[199 : 160] = dep_chan_data_7_31;
    assign token_in_vec_31[4] = token_7_31;
    assign in_chan_dep_vld_vec_31[5] = dep_chan_vld_8_31;
    assign in_chan_dep_data_vec_31[239 : 200] = dep_chan_data_8_31;
    assign token_in_vec_31[5] = token_8_31;
    assign in_chan_dep_vld_vec_31[6] = dep_chan_vld_9_31;
    assign in_chan_dep_data_vec_31[279 : 240] = dep_chan_data_9_31;
    assign token_in_vec_31[6] = token_9_31;
    assign in_chan_dep_vld_vec_31[7] = dep_chan_vld_10_31;
    assign in_chan_dep_data_vec_31[319 : 280] = dep_chan_data_10_31;
    assign token_in_vec_31[7] = token_10_31;
    assign in_chan_dep_vld_vec_31[8] = dep_chan_vld_11_31;
    assign in_chan_dep_data_vec_31[359 : 320] = dep_chan_data_11_31;
    assign token_in_vec_31[8] = token_11_31;
    assign in_chan_dep_vld_vec_31[9] = dep_chan_vld_12_31;
    assign in_chan_dep_data_vec_31[399 : 360] = dep_chan_data_12_31;
    assign token_in_vec_31[9] = token_12_31;
    assign in_chan_dep_vld_vec_31[10] = dep_chan_vld_13_31;
    assign in_chan_dep_data_vec_31[439 : 400] = dep_chan_data_13_31;
    assign token_in_vec_31[10] = token_13_31;
    assign in_chan_dep_vld_vec_31[11] = dep_chan_vld_14_31;
    assign in_chan_dep_data_vec_31[479 : 440] = dep_chan_data_14_31;
    assign token_in_vec_31[11] = token_14_31;
    assign in_chan_dep_vld_vec_31[12] = dep_chan_vld_15_31;
    assign in_chan_dep_data_vec_31[519 : 480] = dep_chan_data_15_31;
    assign token_in_vec_31[12] = token_15_31;
    assign in_chan_dep_vld_vec_31[13] = dep_chan_vld_16_31;
    assign in_chan_dep_data_vec_31[559 : 520] = dep_chan_data_16_31;
    assign token_in_vec_31[13] = token_16_31;
    assign in_chan_dep_vld_vec_31[14] = dep_chan_vld_17_31;
    assign in_chan_dep_data_vec_31[599 : 560] = dep_chan_data_17_31;
    assign token_in_vec_31[14] = token_17_31;
    assign in_chan_dep_vld_vec_31[15] = dep_chan_vld_18_31;
    assign in_chan_dep_data_vec_31[639 : 600] = dep_chan_data_18_31;
    assign token_in_vec_31[15] = token_18_31;
    assign in_chan_dep_vld_vec_31[16] = dep_chan_vld_19_31;
    assign in_chan_dep_data_vec_31[679 : 640] = dep_chan_data_19_31;
    assign token_in_vec_31[16] = token_19_31;
    assign in_chan_dep_vld_vec_31[17] = dep_chan_vld_20_31;
    assign in_chan_dep_data_vec_31[719 : 680] = dep_chan_data_20_31;
    assign token_in_vec_31[17] = token_20_31;
    assign in_chan_dep_vld_vec_31[18] = dep_chan_vld_21_31;
    assign in_chan_dep_data_vec_31[759 : 720] = dep_chan_data_21_31;
    assign token_in_vec_31[18] = token_21_31;
    assign in_chan_dep_vld_vec_31[19] = dep_chan_vld_22_31;
    assign in_chan_dep_data_vec_31[799 : 760] = dep_chan_data_22_31;
    assign token_in_vec_31[19] = token_22_31;
    assign in_chan_dep_vld_vec_31[20] = dep_chan_vld_23_31;
    assign in_chan_dep_data_vec_31[839 : 800] = dep_chan_data_23_31;
    assign token_in_vec_31[20] = token_23_31;
    assign in_chan_dep_vld_vec_31[21] = dep_chan_vld_24_31;
    assign in_chan_dep_data_vec_31[879 : 840] = dep_chan_data_24_31;
    assign token_in_vec_31[21] = token_24_31;
    assign in_chan_dep_vld_vec_31[22] = dep_chan_vld_25_31;
    assign in_chan_dep_data_vec_31[919 : 880] = dep_chan_data_25_31;
    assign token_in_vec_31[22] = token_25_31;
    assign in_chan_dep_vld_vec_31[23] = dep_chan_vld_26_31;
    assign in_chan_dep_data_vec_31[959 : 920] = dep_chan_data_26_31;
    assign token_in_vec_31[23] = token_26_31;
    assign in_chan_dep_vld_vec_31[24] = dep_chan_vld_27_31;
    assign in_chan_dep_data_vec_31[999 : 960] = dep_chan_data_27_31;
    assign token_in_vec_31[24] = token_27_31;
    assign in_chan_dep_vld_vec_31[25] = dep_chan_vld_28_31;
    assign in_chan_dep_data_vec_31[1039 : 1000] = dep_chan_data_28_31;
    assign token_in_vec_31[25] = token_28_31;
    assign in_chan_dep_vld_vec_31[26] = dep_chan_vld_29_31;
    assign in_chan_dep_data_vec_31[1079 : 1040] = dep_chan_data_29_31;
    assign token_in_vec_31[26] = token_29_31;
    assign in_chan_dep_vld_vec_31[27] = dep_chan_vld_30_31;
    assign in_chan_dep_data_vec_31[1119 : 1080] = dep_chan_data_30_31;
    assign token_in_vec_31[27] = token_30_31;
    assign in_chan_dep_vld_vec_31[28] = dep_chan_vld_32_31;
    assign in_chan_dep_data_vec_31[1159 : 1120] = dep_chan_data_32_31;
    assign token_in_vec_31[28] = token_32_31;
    assign in_chan_dep_vld_vec_31[29] = dep_chan_vld_33_31;
    assign in_chan_dep_data_vec_31[1199 : 1160] = dep_chan_data_33_31;
    assign token_in_vec_31[29] = token_33_31;
    assign in_chan_dep_vld_vec_31[30] = dep_chan_vld_34_31;
    assign in_chan_dep_data_vec_31[1239 : 1200] = dep_chan_data_34_31;
    assign token_in_vec_31[30] = token_34_31;
    assign in_chan_dep_vld_vec_31[31] = dep_chan_vld_35_31;
    assign in_chan_dep_data_vec_31[1279 : 1240] = dep_chan_data_35_31;
    assign token_in_vec_31[31] = token_35_31;
    assign in_chan_dep_vld_vec_31[32] = dep_chan_vld_36_31;
    assign in_chan_dep_data_vec_31[1319 : 1280] = dep_chan_data_36_31;
    assign token_in_vec_31[32] = token_36_31;
    assign dep_chan_vld_31_30 = out_chan_dep_vld_vec_31[0];
    assign dep_chan_data_31_30 = out_chan_dep_data_31;
    assign token_31_30 = token_out_vec_31[0];
    assign dep_chan_vld_31_32 = out_chan_dep_vld_vec_31[1];
    assign dep_chan_data_31_32 = out_chan_dep_data_31;
    assign token_31_32 = token_out_vec_31[1];
    assign dep_chan_vld_31_0 = out_chan_dep_vld_vec_31[2];
    assign dep_chan_data_31_0 = out_chan_dep_data_31;
    assign token_31_0 = token_out_vec_31[2];
    assign dep_chan_vld_31_1 = out_chan_dep_vld_vec_31[3];
    assign dep_chan_data_31_1 = out_chan_dep_data_31;
    assign token_31_1 = token_out_vec_31[3];
    assign dep_chan_vld_31_3 = out_chan_dep_vld_vec_31[4];
    assign dep_chan_data_31_3 = out_chan_dep_data_31;
    assign token_31_3 = token_out_vec_31[4];
    assign dep_chan_vld_31_6 = out_chan_dep_vld_vec_31[5];
    assign dep_chan_data_31_6 = out_chan_dep_data_31;
    assign token_31_6 = token_out_vec_31[5];
    assign dep_chan_vld_31_7 = out_chan_dep_vld_vec_31[6];
    assign dep_chan_data_31_7 = out_chan_dep_data_31;
    assign token_31_7 = token_out_vec_31[6];
    assign dep_chan_vld_31_8 = out_chan_dep_vld_vec_31[7];
    assign dep_chan_data_31_8 = out_chan_dep_data_31;
    assign token_31_8 = token_out_vec_31[7];
    assign dep_chan_vld_31_9 = out_chan_dep_vld_vec_31[8];
    assign dep_chan_data_31_9 = out_chan_dep_data_31;
    assign token_31_9 = token_out_vec_31[8];
    assign dep_chan_vld_31_10 = out_chan_dep_vld_vec_31[9];
    assign dep_chan_data_31_10 = out_chan_dep_data_31;
    assign token_31_10 = token_out_vec_31[9];
    assign dep_chan_vld_31_11 = out_chan_dep_vld_vec_31[10];
    assign dep_chan_data_31_11 = out_chan_dep_data_31;
    assign token_31_11 = token_out_vec_31[10];
    assign dep_chan_vld_31_12 = out_chan_dep_vld_vec_31[11];
    assign dep_chan_data_31_12 = out_chan_dep_data_31;
    assign token_31_12 = token_out_vec_31[11];
    assign dep_chan_vld_31_13 = out_chan_dep_vld_vec_31[12];
    assign dep_chan_data_31_13 = out_chan_dep_data_31;
    assign token_31_13 = token_out_vec_31[12];
    assign dep_chan_vld_31_14 = out_chan_dep_vld_vec_31[13];
    assign dep_chan_data_31_14 = out_chan_dep_data_31;
    assign token_31_14 = token_out_vec_31[13];
    assign dep_chan_vld_31_15 = out_chan_dep_vld_vec_31[14];
    assign dep_chan_data_31_15 = out_chan_dep_data_31;
    assign token_31_15 = token_out_vec_31[14];
    assign dep_chan_vld_31_16 = out_chan_dep_vld_vec_31[15];
    assign dep_chan_data_31_16 = out_chan_dep_data_31;
    assign token_31_16 = token_out_vec_31[15];
    assign dep_chan_vld_31_17 = out_chan_dep_vld_vec_31[16];
    assign dep_chan_data_31_17 = out_chan_dep_data_31;
    assign token_31_17 = token_out_vec_31[16];
    assign dep_chan_vld_31_18 = out_chan_dep_vld_vec_31[17];
    assign dep_chan_data_31_18 = out_chan_dep_data_31;
    assign token_31_18 = token_out_vec_31[17];
    assign dep_chan_vld_31_19 = out_chan_dep_vld_vec_31[18];
    assign dep_chan_data_31_19 = out_chan_dep_data_31;
    assign token_31_19 = token_out_vec_31[18];
    assign dep_chan_vld_31_20 = out_chan_dep_vld_vec_31[19];
    assign dep_chan_data_31_20 = out_chan_dep_data_31;
    assign token_31_20 = token_out_vec_31[19];
    assign dep_chan_vld_31_21 = out_chan_dep_vld_vec_31[20];
    assign dep_chan_data_31_21 = out_chan_dep_data_31;
    assign token_31_21 = token_out_vec_31[20];
    assign dep_chan_vld_31_22 = out_chan_dep_vld_vec_31[21];
    assign dep_chan_data_31_22 = out_chan_dep_data_31;
    assign token_31_22 = token_out_vec_31[21];
    assign dep_chan_vld_31_23 = out_chan_dep_vld_vec_31[22];
    assign dep_chan_data_31_23 = out_chan_dep_data_31;
    assign token_31_23 = token_out_vec_31[22];
    assign dep_chan_vld_31_24 = out_chan_dep_vld_vec_31[23];
    assign dep_chan_data_31_24 = out_chan_dep_data_31;
    assign token_31_24 = token_out_vec_31[23];
    assign dep_chan_vld_31_25 = out_chan_dep_vld_vec_31[24];
    assign dep_chan_data_31_25 = out_chan_dep_data_31;
    assign token_31_25 = token_out_vec_31[24];
    assign dep_chan_vld_31_26 = out_chan_dep_vld_vec_31[25];
    assign dep_chan_data_31_26 = out_chan_dep_data_31;
    assign token_31_26 = token_out_vec_31[25];
    assign dep_chan_vld_31_27 = out_chan_dep_vld_vec_31[26];
    assign dep_chan_data_31_27 = out_chan_dep_data_31;
    assign token_31_27 = token_out_vec_31[26];
    assign dep_chan_vld_31_28 = out_chan_dep_vld_vec_31[27];
    assign dep_chan_data_31_28 = out_chan_dep_data_31;
    assign token_31_28 = token_out_vec_31[27];
    assign dep_chan_vld_31_29 = out_chan_dep_vld_vec_31[28];
    assign dep_chan_data_31_29 = out_chan_dep_data_31;
    assign token_31_29 = token_out_vec_31[28];
    assign dep_chan_vld_31_33 = out_chan_dep_vld_vec_31[29];
    assign dep_chan_data_31_33 = out_chan_dep_data_31;
    assign token_31_33 = token_out_vec_31[29];
    assign dep_chan_vld_31_34 = out_chan_dep_vld_vec_31[30];
    assign dep_chan_data_31_34 = out_chan_dep_data_31;
    assign token_31_34 = token_out_vec_31[30];
    assign dep_chan_vld_31_35 = out_chan_dep_vld_vec_31[31];
    assign dep_chan_data_31_35 = out_chan_dep_data_31;
    assign token_31_35 = token_out_vec_31[31];
    assign dep_chan_vld_31_36 = out_chan_dep_vld_vec_31[32];
    assign dep_chan_data_31_36 = out_chan_dep_data_31;
    assign token_31_36 = token_out_vec_31[32];

    // Process: ProcessingElement_27_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 32, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_32 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_32),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_32),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_32),
        .token_in_vec(token_in_vec_32),
        .dl_detect_in(dl_detect_out),
        .origin(origin[32]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_32),
        .out_chan_dep_data(out_chan_dep_data_32),
        .token_out_vec(token_out_vec_32),
        .dl_detect_out(dl_in_vec[32]));

    assign proc_32_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_26_blk_n) | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_26_blk_n) | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_WriteC_Flattened_fu_179.cPipes_26_blk_n);
    assign proc_32_data_PIPO_blk[0] = 1'b0;
    assign proc_32_start_FIFO_blk[0] = 1'b0;
    assign proc_32_TLF_FIFO_blk[0] = 1'b0;
    assign proc_32_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_32_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_32[0] = dl_detect_out ? proc_dep_vld_vec_32_reg[0] : (proc_32_data_FIFO_blk[0] | proc_32_data_PIPO_blk[0] | proc_32_start_FIFO_blk[0] | proc_32_TLF_FIFO_blk[0] | proc_32_input_sync_blk[0] | proc_32_output_sync_blk[0]);
    assign proc_32_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_27_blk_n) | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_27_blk_n) | (~ProcessingElement_27_U0.grp_ProcessingElement_27_Pipeline_WriteC_Flattened_fu_179.cPipes_27_blk_n);
    assign proc_32_data_PIPO_blk[1] = 1'b0;
    assign proc_32_start_FIFO_blk[1] = 1'b0;
    assign proc_32_TLF_FIFO_blk[1] = 1'b0;
    assign proc_32_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_32_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_32[1] = dl_detect_out ? proc_dep_vld_vec_32_reg[1] : (proc_32_data_FIFO_blk[1] | proc_32_data_PIPO_blk[1] | proc_32_start_FIFO_blk[1] | proc_32_TLF_FIFO_blk[1] | proc_32_input_sync_blk[1] | proc_32_output_sync_blk[1]);
    assign proc_32_data_FIFO_blk[2] = 1'b0;
    assign proc_32_data_PIPO_blk[2] = 1'b0;
    assign proc_32_start_FIFO_blk[2] = 1'b0;
    assign proc_32_TLF_FIFO_blk[2] = 1'b0;
    assign proc_32_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_32_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_32[2] = dl_detect_out ? proc_dep_vld_vec_32_reg[2] : (proc_32_data_FIFO_blk[2] | proc_32_data_PIPO_blk[2] | proc_32_start_FIFO_blk[2] | proc_32_TLF_FIFO_blk[2] | proc_32_input_sync_blk[2] | proc_32_output_sync_blk[2]);
    assign proc_32_data_FIFO_blk[3] = 1'b0;
    assign proc_32_data_PIPO_blk[3] = 1'b0;
    assign proc_32_start_FIFO_blk[3] = 1'b0;
    assign proc_32_TLF_FIFO_blk[3] = 1'b0;
    assign proc_32_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_32_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_32[3] = dl_detect_out ? proc_dep_vld_vec_32_reg[3] : (proc_32_data_FIFO_blk[3] | proc_32_data_PIPO_blk[3] | proc_32_start_FIFO_blk[3] | proc_32_TLF_FIFO_blk[3] | proc_32_input_sync_blk[3] | proc_32_output_sync_blk[3]);
    assign proc_32_data_FIFO_blk[4] = 1'b0;
    assign proc_32_data_PIPO_blk[4] = 1'b0;
    assign proc_32_start_FIFO_blk[4] = 1'b0;
    assign proc_32_TLF_FIFO_blk[4] = 1'b0;
    assign proc_32_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_32_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_32[4] = dl_detect_out ? proc_dep_vld_vec_32_reg[4] : (proc_32_data_FIFO_blk[4] | proc_32_data_PIPO_blk[4] | proc_32_start_FIFO_blk[4] | proc_32_TLF_FIFO_blk[4] | proc_32_input_sync_blk[4] | proc_32_output_sync_blk[4]);
    assign proc_32_data_FIFO_blk[5] = 1'b0;
    assign proc_32_data_PIPO_blk[5] = 1'b0;
    assign proc_32_start_FIFO_blk[5] = 1'b0;
    assign proc_32_TLF_FIFO_blk[5] = 1'b0;
    assign proc_32_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_32_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_32[5] = dl_detect_out ? proc_dep_vld_vec_32_reg[5] : (proc_32_data_FIFO_blk[5] | proc_32_data_PIPO_blk[5] | proc_32_start_FIFO_blk[5] | proc_32_TLF_FIFO_blk[5] | proc_32_input_sync_blk[5] | proc_32_output_sync_blk[5]);
    assign proc_32_data_FIFO_blk[6] = 1'b0;
    assign proc_32_data_PIPO_blk[6] = 1'b0;
    assign proc_32_start_FIFO_blk[6] = 1'b0;
    assign proc_32_TLF_FIFO_blk[6] = 1'b0;
    assign proc_32_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_32_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_32[6] = dl_detect_out ? proc_dep_vld_vec_32_reg[6] : (proc_32_data_FIFO_blk[6] | proc_32_data_PIPO_blk[6] | proc_32_start_FIFO_blk[6] | proc_32_TLF_FIFO_blk[6] | proc_32_input_sync_blk[6] | proc_32_output_sync_blk[6]);
    assign proc_32_data_FIFO_blk[7] = 1'b0;
    assign proc_32_data_PIPO_blk[7] = 1'b0;
    assign proc_32_start_FIFO_blk[7] = 1'b0;
    assign proc_32_TLF_FIFO_blk[7] = 1'b0;
    assign proc_32_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_32_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_32[7] = dl_detect_out ? proc_dep_vld_vec_32_reg[7] : (proc_32_data_FIFO_blk[7] | proc_32_data_PIPO_blk[7] | proc_32_start_FIFO_blk[7] | proc_32_TLF_FIFO_blk[7] | proc_32_input_sync_blk[7] | proc_32_output_sync_blk[7]);
    assign proc_32_data_FIFO_blk[8] = 1'b0;
    assign proc_32_data_PIPO_blk[8] = 1'b0;
    assign proc_32_start_FIFO_blk[8] = 1'b0;
    assign proc_32_TLF_FIFO_blk[8] = 1'b0;
    assign proc_32_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_32_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_32[8] = dl_detect_out ? proc_dep_vld_vec_32_reg[8] : (proc_32_data_FIFO_blk[8] | proc_32_data_PIPO_blk[8] | proc_32_start_FIFO_blk[8] | proc_32_TLF_FIFO_blk[8] | proc_32_input_sync_blk[8] | proc_32_output_sync_blk[8]);
    assign proc_32_data_FIFO_blk[9] = 1'b0;
    assign proc_32_data_PIPO_blk[9] = 1'b0;
    assign proc_32_start_FIFO_blk[9] = 1'b0;
    assign proc_32_TLF_FIFO_blk[9] = 1'b0;
    assign proc_32_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_32_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_32[9] = dl_detect_out ? proc_dep_vld_vec_32_reg[9] : (proc_32_data_FIFO_blk[9] | proc_32_data_PIPO_blk[9] | proc_32_start_FIFO_blk[9] | proc_32_TLF_FIFO_blk[9] | proc_32_input_sync_blk[9] | proc_32_output_sync_blk[9]);
    assign proc_32_data_FIFO_blk[10] = 1'b0;
    assign proc_32_data_PIPO_blk[10] = 1'b0;
    assign proc_32_start_FIFO_blk[10] = 1'b0;
    assign proc_32_TLF_FIFO_blk[10] = 1'b0;
    assign proc_32_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_32_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_32[10] = dl_detect_out ? proc_dep_vld_vec_32_reg[10] : (proc_32_data_FIFO_blk[10] | proc_32_data_PIPO_blk[10] | proc_32_start_FIFO_blk[10] | proc_32_TLF_FIFO_blk[10] | proc_32_input_sync_blk[10] | proc_32_output_sync_blk[10]);
    assign proc_32_data_FIFO_blk[11] = 1'b0;
    assign proc_32_data_PIPO_blk[11] = 1'b0;
    assign proc_32_start_FIFO_blk[11] = 1'b0;
    assign proc_32_TLF_FIFO_blk[11] = 1'b0;
    assign proc_32_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_32_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_32[11] = dl_detect_out ? proc_dep_vld_vec_32_reg[11] : (proc_32_data_FIFO_blk[11] | proc_32_data_PIPO_blk[11] | proc_32_start_FIFO_blk[11] | proc_32_TLF_FIFO_blk[11] | proc_32_input_sync_blk[11] | proc_32_output_sync_blk[11]);
    assign proc_32_data_FIFO_blk[12] = 1'b0;
    assign proc_32_data_PIPO_blk[12] = 1'b0;
    assign proc_32_start_FIFO_blk[12] = 1'b0;
    assign proc_32_TLF_FIFO_blk[12] = 1'b0;
    assign proc_32_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_32_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_32[12] = dl_detect_out ? proc_dep_vld_vec_32_reg[12] : (proc_32_data_FIFO_blk[12] | proc_32_data_PIPO_blk[12] | proc_32_start_FIFO_blk[12] | proc_32_TLF_FIFO_blk[12] | proc_32_input_sync_blk[12] | proc_32_output_sync_blk[12]);
    assign proc_32_data_FIFO_blk[13] = 1'b0;
    assign proc_32_data_PIPO_blk[13] = 1'b0;
    assign proc_32_start_FIFO_blk[13] = 1'b0;
    assign proc_32_TLF_FIFO_blk[13] = 1'b0;
    assign proc_32_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_32_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_32[13] = dl_detect_out ? proc_dep_vld_vec_32_reg[13] : (proc_32_data_FIFO_blk[13] | proc_32_data_PIPO_blk[13] | proc_32_start_FIFO_blk[13] | proc_32_TLF_FIFO_blk[13] | proc_32_input_sync_blk[13] | proc_32_output_sync_blk[13]);
    assign proc_32_data_FIFO_blk[14] = 1'b0;
    assign proc_32_data_PIPO_blk[14] = 1'b0;
    assign proc_32_start_FIFO_blk[14] = 1'b0;
    assign proc_32_TLF_FIFO_blk[14] = 1'b0;
    assign proc_32_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_32_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_32[14] = dl_detect_out ? proc_dep_vld_vec_32_reg[14] : (proc_32_data_FIFO_blk[14] | proc_32_data_PIPO_blk[14] | proc_32_start_FIFO_blk[14] | proc_32_TLF_FIFO_blk[14] | proc_32_input_sync_blk[14] | proc_32_output_sync_blk[14]);
    assign proc_32_data_FIFO_blk[15] = 1'b0;
    assign proc_32_data_PIPO_blk[15] = 1'b0;
    assign proc_32_start_FIFO_blk[15] = 1'b0;
    assign proc_32_TLF_FIFO_blk[15] = 1'b0;
    assign proc_32_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_32_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_32[15] = dl_detect_out ? proc_dep_vld_vec_32_reg[15] : (proc_32_data_FIFO_blk[15] | proc_32_data_PIPO_blk[15] | proc_32_start_FIFO_blk[15] | proc_32_TLF_FIFO_blk[15] | proc_32_input_sync_blk[15] | proc_32_output_sync_blk[15]);
    assign proc_32_data_FIFO_blk[16] = 1'b0;
    assign proc_32_data_PIPO_blk[16] = 1'b0;
    assign proc_32_start_FIFO_blk[16] = 1'b0;
    assign proc_32_TLF_FIFO_blk[16] = 1'b0;
    assign proc_32_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_32_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_32[16] = dl_detect_out ? proc_dep_vld_vec_32_reg[16] : (proc_32_data_FIFO_blk[16] | proc_32_data_PIPO_blk[16] | proc_32_start_FIFO_blk[16] | proc_32_TLF_FIFO_blk[16] | proc_32_input_sync_blk[16] | proc_32_output_sync_blk[16]);
    assign proc_32_data_FIFO_blk[17] = 1'b0;
    assign proc_32_data_PIPO_blk[17] = 1'b0;
    assign proc_32_start_FIFO_blk[17] = 1'b0;
    assign proc_32_TLF_FIFO_blk[17] = 1'b0;
    assign proc_32_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_32_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_32[17] = dl_detect_out ? proc_dep_vld_vec_32_reg[17] : (proc_32_data_FIFO_blk[17] | proc_32_data_PIPO_blk[17] | proc_32_start_FIFO_blk[17] | proc_32_TLF_FIFO_blk[17] | proc_32_input_sync_blk[17] | proc_32_output_sync_blk[17]);
    assign proc_32_data_FIFO_blk[18] = 1'b0;
    assign proc_32_data_PIPO_blk[18] = 1'b0;
    assign proc_32_start_FIFO_blk[18] = 1'b0;
    assign proc_32_TLF_FIFO_blk[18] = 1'b0;
    assign proc_32_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_32_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_32[18] = dl_detect_out ? proc_dep_vld_vec_32_reg[18] : (proc_32_data_FIFO_blk[18] | proc_32_data_PIPO_blk[18] | proc_32_start_FIFO_blk[18] | proc_32_TLF_FIFO_blk[18] | proc_32_input_sync_blk[18] | proc_32_output_sync_blk[18]);
    assign proc_32_data_FIFO_blk[19] = 1'b0;
    assign proc_32_data_PIPO_blk[19] = 1'b0;
    assign proc_32_start_FIFO_blk[19] = 1'b0;
    assign proc_32_TLF_FIFO_blk[19] = 1'b0;
    assign proc_32_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_32_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_32[19] = dl_detect_out ? proc_dep_vld_vec_32_reg[19] : (proc_32_data_FIFO_blk[19] | proc_32_data_PIPO_blk[19] | proc_32_start_FIFO_blk[19] | proc_32_TLF_FIFO_blk[19] | proc_32_input_sync_blk[19] | proc_32_output_sync_blk[19]);
    assign proc_32_data_FIFO_blk[20] = 1'b0;
    assign proc_32_data_PIPO_blk[20] = 1'b0;
    assign proc_32_start_FIFO_blk[20] = 1'b0;
    assign proc_32_TLF_FIFO_blk[20] = 1'b0;
    assign proc_32_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_32_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_32[20] = dl_detect_out ? proc_dep_vld_vec_32_reg[20] : (proc_32_data_FIFO_blk[20] | proc_32_data_PIPO_blk[20] | proc_32_start_FIFO_blk[20] | proc_32_TLF_FIFO_blk[20] | proc_32_input_sync_blk[20] | proc_32_output_sync_blk[20]);
    assign proc_32_data_FIFO_blk[21] = 1'b0;
    assign proc_32_data_PIPO_blk[21] = 1'b0;
    assign proc_32_start_FIFO_blk[21] = 1'b0;
    assign proc_32_TLF_FIFO_blk[21] = 1'b0;
    assign proc_32_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_32_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_32[21] = dl_detect_out ? proc_dep_vld_vec_32_reg[21] : (proc_32_data_FIFO_blk[21] | proc_32_data_PIPO_blk[21] | proc_32_start_FIFO_blk[21] | proc_32_TLF_FIFO_blk[21] | proc_32_input_sync_blk[21] | proc_32_output_sync_blk[21]);
    assign proc_32_data_FIFO_blk[22] = 1'b0;
    assign proc_32_data_PIPO_blk[22] = 1'b0;
    assign proc_32_start_FIFO_blk[22] = 1'b0;
    assign proc_32_TLF_FIFO_blk[22] = 1'b0;
    assign proc_32_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_32_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_32[22] = dl_detect_out ? proc_dep_vld_vec_32_reg[22] : (proc_32_data_FIFO_blk[22] | proc_32_data_PIPO_blk[22] | proc_32_start_FIFO_blk[22] | proc_32_TLF_FIFO_blk[22] | proc_32_input_sync_blk[22] | proc_32_output_sync_blk[22]);
    assign proc_32_data_FIFO_blk[23] = 1'b0;
    assign proc_32_data_PIPO_blk[23] = 1'b0;
    assign proc_32_start_FIFO_blk[23] = 1'b0;
    assign proc_32_TLF_FIFO_blk[23] = 1'b0;
    assign proc_32_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_32_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_32[23] = dl_detect_out ? proc_dep_vld_vec_32_reg[23] : (proc_32_data_FIFO_blk[23] | proc_32_data_PIPO_blk[23] | proc_32_start_FIFO_blk[23] | proc_32_TLF_FIFO_blk[23] | proc_32_input_sync_blk[23] | proc_32_output_sync_blk[23]);
    assign proc_32_data_FIFO_blk[24] = 1'b0;
    assign proc_32_data_PIPO_blk[24] = 1'b0;
    assign proc_32_start_FIFO_blk[24] = 1'b0;
    assign proc_32_TLF_FIFO_blk[24] = 1'b0;
    assign proc_32_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_32_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_32[24] = dl_detect_out ? proc_dep_vld_vec_32_reg[24] : (proc_32_data_FIFO_blk[24] | proc_32_data_PIPO_blk[24] | proc_32_start_FIFO_blk[24] | proc_32_TLF_FIFO_blk[24] | proc_32_input_sync_blk[24] | proc_32_output_sync_blk[24]);
    assign proc_32_data_FIFO_blk[25] = 1'b0;
    assign proc_32_data_PIPO_blk[25] = 1'b0;
    assign proc_32_start_FIFO_blk[25] = 1'b0;
    assign proc_32_TLF_FIFO_blk[25] = 1'b0;
    assign proc_32_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_32_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_32[25] = dl_detect_out ? proc_dep_vld_vec_32_reg[25] : (proc_32_data_FIFO_blk[25] | proc_32_data_PIPO_blk[25] | proc_32_start_FIFO_blk[25] | proc_32_TLF_FIFO_blk[25] | proc_32_input_sync_blk[25] | proc_32_output_sync_blk[25]);
    assign proc_32_data_FIFO_blk[26] = 1'b0;
    assign proc_32_data_PIPO_blk[26] = 1'b0;
    assign proc_32_start_FIFO_blk[26] = 1'b0;
    assign proc_32_TLF_FIFO_blk[26] = 1'b0;
    assign proc_32_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_32_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_32[26] = dl_detect_out ? proc_dep_vld_vec_32_reg[26] : (proc_32_data_FIFO_blk[26] | proc_32_data_PIPO_blk[26] | proc_32_start_FIFO_blk[26] | proc_32_TLF_FIFO_blk[26] | proc_32_input_sync_blk[26] | proc_32_output_sync_blk[26]);
    assign proc_32_data_FIFO_blk[27] = 1'b0;
    assign proc_32_data_PIPO_blk[27] = 1'b0;
    assign proc_32_start_FIFO_blk[27] = 1'b0;
    assign proc_32_TLF_FIFO_blk[27] = 1'b0;
    assign proc_32_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_32_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_32[27] = dl_detect_out ? proc_dep_vld_vec_32_reg[27] : (proc_32_data_FIFO_blk[27] | proc_32_data_PIPO_blk[27] | proc_32_start_FIFO_blk[27] | proc_32_TLF_FIFO_blk[27] | proc_32_input_sync_blk[27] | proc_32_output_sync_blk[27]);
    assign proc_32_data_FIFO_blk[28] = 1'b0;
    assign proc_32_data_PIPO_blk[28] = 1'b0;
    assign proc_32_start_FIFO_blk[28] = 1'b0;
    assign proc_32_TLF_FIFO_blk[28] = 1'b0;
    assign proc_32_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_32_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_32[28] = dl_detect_out ? proc_dep_vld_vec_32_reg[28] : (proc_32_data_FIFO_blk[28] | proc_32_data_PIPO_blk[28] | proc_32_start_FIFO_blk[28] | proc_32_TLF_FIFO_blk[28] | proc_32_input_sync_blk[28] | proc_32_output_sync_blk[28]);
    assign proc_32_data_FIFO_blk[29] = 1'b0;
    assign proc_32_data_PIPO_blk[29] = 1'b0;
    assign proc_32_start_FIFO_blk[29] = 1'b0;
    assign proc_32_TLF_FIFO_blk[29] = 1'b0;
    assign proc_32_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_32_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_32[29] = dl_detect_out ? proc_dep_vld_vec_32_reg[29] : (proc_32_data_FIFO_blk[29] | proc_32_data_PIPO_blk[29] | proc_32_start_FIFO_blk[29] | proc_32_TLF_FIFO_blk[29] | proc_32_input_sync_blk[29] | proc_32_output_sync_blk[29]);
    assign proc_32_data_FIFO_blk[30] = 1'b0;
    assign proc_32_data_PIPO_blk[30] = 1'b0;
    assign proc_32_start_FIFO_blk[30] = 1'b0;
    assign proc_32_TLF_FIFO_blk[30] = 1'b0;
    assign proc_32_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_32_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_32[30] = dl_detect_out ? proc_dep_vld_vec_32_reg[30] : (proc_32_data_FIFO_blk[30] | proc_32_data_PIPO_blk[30] | proc_32_start_FIFO_blk[30] | proc_32_TLF_FIFO_blk[30] | proc_32_input_sync_blk[30] | proc_32_output_sync_blk[30]);
    assign proc_32_data_FIFO_blk[31] = 1'b0;
    assign proc_32_data_PIPO_blk[31] = 1'b0;
    assign proc_32_start_FIFO_blk[31] = 1'b0;
    assign proc_32_TLF_FIFO_blk[31] = 1'b0;
    assign proc_32_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_32_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_32[31] = dl_detect_out ? proc_dep_vld_vec_32_reg[31] : (proc_32_data_FIFO_blk[31] | proc_32_data_PIPO_blk[31] | proc_32_start_FIFO_blk[31] | proc_32_TLF_FIFO_blk[31] | proc_32_input_sync_blk[31] | proc_32_output_sync_blk[31]);
    assign proc_32_data_FIFO_blk[32] = 1'b0;
    assign proc_32_data_PIPO_blk[32] = 1'b0;
    assign proc_32_start_FIFO_blk[32] = 1'b0;
    assign proc_32_TLF_FIFO_blk[32] = 1'b0;
    assign proc_32_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_27_U0_ap_ready & ProcessingElement_27_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_32_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_32[32] = dl_detect_out ? proc_dep_vld_vec_32_reg[32] : (proc_32_data_FIFO_blk[32] | proc_32_data_PIPO_blk[32] | proc_32_start_FIFO_blk[32] | proc_32_TLF_FIFO_blk[32] | proc_32_input_sync_blk[32] | proc_32_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_32_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_32_reg <= proc_dep_vld_vec_32;
        end
    end
    assign in_chan_dep_vld_vec_32[0] = dep_chan_vld_0_32;
    assign in_chan_dep_data_vec_32[39 : 0] = dep_chan_data_0_32;
    assign token_in_vec_32[0] = token_0_32;
    assign in_chan_dep_vld_vec_32[1] = dep_chan_vld_1_32;
    assign in_chan_dep_data_vec_32[79 : 40] = dep_chan_data_1_32;
    assign token_in_vec_32[1] = token_1_32;
    assign in_chan_dep_vld_vec_32[2] = dep_chan_vld_3_32;
    assign in_chan_dep_data_vec_32[119 : 80] = dep_chan_data_3_32;
    assign token_in_vec_32[2] = token_3_32;
    assign in_chan_dep_vld_vec_32[3] = dep_chan_vld_6_32;
    assign in_chan_dep_data_vec_32[159 : 120] = dep_chan_data_6_32;
    assign token_in_vec_32[3] = token_6_32;
    assign in_chan_dep_vld_vec_32[4] = dep_chan_vld_7_32;
    assign in_chan_dep_data_vec_32[199 : 160] = dep_chan_data_7_32;
    assign token_in_vec_32[4] = token_7_32;
    assign in_chan_dep_vld_vec_32[5] = dep_chan_vld_8_32;
    assign in_chan_dep_data_vec_32[239 : 200] = dep_chan_data_8_32;
    assign token_in_vec_32[5] = token_8_32;
    assign in_chan_dep_vld_vec_32[6] = dep_chan_vld_9_32;
    assign in_chan_dep_data_vec_32[279 : 240] = dep_chan_data_9_32;
    assign token_in_vec_32[6] = token_9_32;
    assign in_chan_dep_vld_vec_32[7] = dep_chan_vld_10_32;
    assign in_chan_dep_data_vec_32[319 : 280] = dep_chan_data_10_32;
    assign token_in_vec_32[7] = token_10_32;
    assign in_chan_dep_vld_vec_32[8] = dep_chan_vld_11_32;
    assign in_chan_dep_data_vec_32[359 : 320] = dep_chan_data_11_32;
    assign token_in_vec_32[8] = token_11_32;
    assign in_chan_dep_vld_vec_32[9] = dep_chan_vld_12_32;
    assign in_chan_dep_data_vec_32[399 : 360] = dep_chan_data_12_32;
    assign token_in_vec_32[9] = token_12_32;
    assign in_chan_dep_vld_vec_32[10] = dep_chan_vld_13_32;
    assign in_chan_dep_data_vec_32[439 : 400] = dep_chan_data_13_32;
    assign token_in_vec_32[10] = token_13_32;
    assign in_chan_dep_vld_vec_32[11] = dep_chan_vld_14_32;
    assign in_chan_dep_data_vec_32[479 : 440] = dep_chan_data_14_32;
    assign token_in_vec_32[11] = token_14_32;
    assign in_chan_dep_vld_vec_32[12] = dep_chan_vld_15_32;
    assign in_chan_dep_data_vec_32[519 : 480] = dep_chan_data_15_32;
    assign token_in_vec_32[12] = token_15_32;
    assign in_chan_dep_vld_vec_32[13] = dep_chan_vld_16_32;
    assign in_chan_dep_data_vec_32[559 : 520] = dep_chan_data_16_32;
    assign token_in_vec_32[13] = token_16_32;
    assign in_chan_dep_vld_vec_32[14] = dep_chan_vld_17_32;
    assign in_chan_dep_data_vec_32[599 : 560] = dep_chan_data_17_32;
    assign token_in_vec_32[14] = token_17_32;
    assign in_chan_dep_vld_vec_32[15] = dep_chan_vld_18_32;
    assign in_chan_dep_data_vec_32[639 : 600] = dep_chan_data_18_32;
    assign token_in_vec_32[15] = token_18_32;
    assign in_chan_dep_vld_vec_32[16] = dep_chan_vld_19_32;
    assign in_chan_dep_data_vec_32[679 : 640] = dep_chan_data_19_32;
    assign token_in_vec_32[16] = token_19_32;
    assign in_chan_dep_vld_vec_32[17] = dep_chan_vld_20_32;
    assign in_chan_dep_data_vec_32[719 : 680] = dep_chan_data_20_32;
    assign token_in_vec_32[17] = token_20_32;
    assign in_chan_dep_vld_vec_32[18] = dep_chan_vld_21_32;
    assign in_chan_dep_data_vec_32[759 : 720] = dep_chan_data_21_32;
    assign token_in_vec_32[18] = token_21_32;
    assign in_chan_dep_vld_vec_32[19] = dep_chan_vld_22_32;
    assign in_chan_dep_data_vec_32[799 : 760] = dep_chan_data_22_32;
    assign token_in_vec_32[19] = token_22_32;
    assign in_chan_dep_vld_vec_32[20] = dep_chan_vld_23_32;
    assign in_chan_dep_data_vec_32[839 : 800] = dep_chan_data_23_32;
    assign token_in_vec_32[20] = token_23_32;
    assign in_chan_dep_vld_vec_32[21] = dep_chan_vld_24_32;
    assign in_chan_dep_data_vec_32[879 : 840] = dep_chan_data_24_32;
    assign token_in_vec_32[21] = token_24_32;
    assign in_chan_dep_vld_vec_32[22] = dep_chan_vld_25_32;
    assign in_chan_dep_data_vec_32[919 : 880] = dep_chan_data_25_32;
    assign token_in_vec_32[22] = token_25_32;
    assign in_chan_dep_vld_vec_32[23] = dep_chan_vld_26_32;
    assign in_chan_dep_data_vec_32[959 : 920] = dep_chan_data_26_32;
    assign token_in_vec_32[23] = token_26_32;
    assign in_chan_dep_vld_vec_32[24] = dep_chan_vld_27_32;
    assign in_chan_dep_data_vec_32[999 : 960] = dep_chan_data_27_32;
    assign token_in_vec_32[24] = token_27_32;
    assign in_chan_dep_vld_vec_32[25] = dep_chan_vld_28_32;
    assign in_chan_dep_data_vec_32[1039 : 1000] = dep_chan_data_28_32;
    assign token_in_vec_32[25] = token_28_32;
    assign in_chan_dep_vld_vec_32[26] = dep_chan_vld_29_32;
    assign in_chan_dep_data_vec_32[1079 : 1040] = dep_chan_data_29_32;
    assign token_in_vec_32[26] = token_29_32;
    assign in_chan_dep_vld_vec_32[27] = dep_chan_vld_30_32;
    assign in_chan_dep_data_vec_32[1119 : 1080] = dep_chan_data_30_32;
    assign token_in_vec_32[27] = token_30_32;
    assign in_chan_dep_vld_vec_32[28] = dep_chan_vld_31_32;
    assign in_chan_dep_data_vec_32[1159 : 1120] = dep_chan_data_31_32;
    assign token_in_vec_32[28] = token_31_32;
    assign in_chan_dep_vld_vec_32[29] = dep_chan_vld_33_32;
    assign in_chan_dep_data_vec_32[1199 : 1160] = dep_chan_data_33_32;
    assign token_in_vec_32[29] = token_33_32;
    assign in_chan_dep_vld_vec_32[30] = dep_chan_vld_34_32;
    assign in_chan_dep_data_vec_32[1239 : 1200] = dep_chan_data_34_32;
    assign token_in_vec_32[30] = token_34_32;
    assign in_chan_dep_vld_vec_32[31] = dep_chan_vld_35_32;
    assign in_chan_dep_data_vec_32[1279 : 1240] = dep_chan_data_35_32;
    assign token_in_vec_32[31] = token_35_32;
    assign in_chan_dep_vld_vec_32[32] = dep_chan_vld_36_32;
    assign in_chan_dep_data_vec_32[1319 : 1280] = dep_chan_data_36_32;
    assign token_in_vec_32[32] = token_36_32;
    assign dep_chan_vld_32_31 = out_chan_dep_vld_vec_32[0];
    assign dep_chan_data_32_31 = out_chan_dep_data_32;
    assign token_32_31 = token_out_vec_32[0];
    assign dep_chan_vld_32_33 = out_chan_dep_vld_vec_32[1];
    assign dep_chan_data_32_33 = out_chan_dep_data_32;
    assign token_32_33 = token_out_vec_32[1];
    assign dep_chan_vld_32_0 = out_chan_dep_vld_vec_32[2];
    assign dep_chan_data_32_0 = out_chan_dep_data_32;
    assign token_32_0 = token_out_vec_32[2];
    assign dep_chan_vld_32_1 = out_chan_dep_vld_vec_32[3];
    assign dep_chan_data_32_1 = out_chan_dep_data_32;
    assign token_32_1 = token_out_vec_32[3];
    assign dep_chan_vld_32_3 = out_chan_dep_vld_vec_32[4];
    assign dep_chan_data_32_3 = out_chan_dep_data_32;
    assign token_32_3 = token_out_vec_32[4];
    assign dep_chan_vld_32_6 = out_chan_dep_vld_vec_32[5];
    assign dep_chan_data_32_6 = out_chan_dep_data_32;
    assign token_32_6 = token_out_vec_32[5];
    assign dep_chan_vld_32_7 = out_chan_dep_vld_vec_32[6];
    assign dep_chan_data_32_7 = out_chan_dep_data_32;
    assign token_32_7 = token_out_vec_32[6];
    assign dep_chan_vld_32_8 = out_chan_dep_vld_vec_32[7];
    assign dep_chan_data_32_8 = out_chan_dep_data_32;
    assign token_32_8 = token_out_vec_32[7];
    assign dep_chan_vld_32_9 = out_chan_dep_vld_vec_32[8];
    assign dep_chan_data_32_9 = out_chan_dep_data_32;
    assign token_32_9 = token_out_vec_32[8];
    assign dep_chan_vld_32_10 = out_chan_dep_vld_vec_32[9];
    assign dep_chan_data_32_10 = out_chan_dep_data_32;
    assign token_32_10 = token_out_vec_32[9];
    assign dep_chan_vld_32_11 = out_chan_dep_vld_vec_32[10];
    assign dep_chan_data_32_11 = out_chan_dep_data_32;
    assign token_32_11 = token_out_vec_32[10];
    assign dep_chan_vld_32_12 = out_chan_dep_vld_vec_32[11];
    assign dep_chan_data_32_12 = out_chan_dep_data_32;
    assign token_32_12 = token_out_vec_32[11];
    assign dep_chan_vld_32_13 = out_chan_dep_vld_vec_32[12];
    assign dep_chan_data_32_13 = out_chan_dep_data_32;
    assign token_32_13 = token_out_vec_32[12];
    assign dep_chan_vld_32_14 = out_chan_dep_vld_vec_32[13];
    assign dep_chan_data_32_14 = out_chan_dep_data_32;
    assign token_32_14 = token_out_vec_32[13];
    assign dep_chan_vld_32_15 = out_chan_dep_vld_vec_32[14];
    assign dep_chan_data_32_15 = out_chan_dep_data_32;
    assign token_32_15 = token_out_vec_32[14];
    assign dep_chan_vld_32_16 = out_chan_dep_vld_vec_32[15];
    assign dep_chan_data_32_16 = out_chan_dep_data_32;
    assign token_32_16 = token_out_vec_32[15];
    assign dep_chan_vld_32_17 = out_chan_dep_vld_vec_32[16];
    assign dep_chan_data_32_17 = out_chan_dep_data_32;
    assign token_32_17 = token_out_vec_32[16];
    assign dep_chan_vld_32_18 = out_chan_dep_vld_vec_32[17];
    assign dep_chan_data_32_18 = out_chan_dep_data_32;
    assign token_32_18 = token_out_vec_32[17];
    assign dep_chan_vld_32_19 = out_chan_dep_vld_vec_32[18];
    assign dep_chan_data_32_19 = out_chan_dep_data_32;
    assign token_32_19 = token_out_vec_32[18];
    assign dep_chan_vld_32_20 = out_chan_dep_vld_vec_32[19];
    assign dep_chan_data_32_20 = out_chan_dep_data_32;
    assign token_32_20 = token_out_vec_32[19];
    assign dep_chan_vld_32_21 = out_chan_dep_vld_vec_32[20];
    assign dep_chan_data_32_21 = out_chan_dep_data_32;
    assign token_32_21 = token_out_vec_32[20];
    assign dep_chan_vld_32_22 = out_chan_dep_vld_vec_32[21];
    assign dep_chan_data_32_22 = out_chan_dep_data_32;
    assign token_32_22 = token_out_vec_32[21];
    assign dep_chan_vld_32_23 = out_chan_dep_vld_vec_32[22];
    assign dep_chan_data_32_23 = out_chan_dep_data_32;
    assign token_32_23 = token_out_vec_32[22];
    assign dep_chan_vld_32_24 = out_chan_dep_vld_vec_32[23];
    assign dep_chan_data_32_24 = out_chan_dep_data_32;
    assign token_32_24 = token_out_vec_32[23];
    assign dep_chan_vld_32_25 = out_chan_dep_vld_vec_32[24];
    assign dep_chan_data_32_25 = out_chan_dep_data_32;
    assign token_32_25 = token_out_vec_32[24];
    assign dep_chan_vld_32_26 = out_chan_dep_vld_vec_32[25];
    assign dep_chan_data_32_26 = out_chan_dep_data_32;
    assign token_32_26 = token_out_vec_32[25];
    assign dep_chan_vld_32_27 = out_chan_dep_vld_vec_32[26];
    assign dep_chan_data_32_27 = out_chan_dep_data_32;
    assign token_32_27 = token_out_vec_32[26];
    assign dep_chan_vld_32_28 = out_chan_dep_vld_vec_32[27];
    assign dep_chan_data_32_28 = out_chan_dep_data_32;
    assign token_32_28 = token_out_vec_32[27];
    assign dep_chan_vld_32_29 = out_chan_dep_vld_vec_32[28];
    assign dep_chan_data_32_29 = out_chan_dep_data_32;
    assign token_32_29 = token_out_vec_32[28];
    assign dep_chan_vld_32_30 = out_chan_dep_vld_vec_32[29];
    assign dep_chan_data_32_30 = out_chan_dep_data_32;
    assign token_32_30 = token_out_vec_32[29];
    assign dep_chan_vld_32_34 = out_chan_dep_vld_vec_32[30];
    assign dep_chan_data_32_34 = out_chan_dep_data_32;
    assign token_32_34 = token_out_vec_32[30];
    assign dep_chan_vld_32_35 = out_chan_dep_vld_vec_32[31];
    assign dep_chan_data_32_35 = out_chan_dep_data_32;
    assign token_32_35 = token_out_vec_32[31];
    assign dep_chan_vld_32_36 = out_chan_dep_vld_vec_32[32];
    assign dep_chan_data_32_36 = out_chan_dep_data_32;
    assign token_32_36 = token_out_vec_32[32];

    // Process: ProcessingElement_28_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 33, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_33 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_33),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_33),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_33),
        .token_in_vec(token_in_vec_33),
        .dl_detect_in(dl_detect_out),
        .origin(origin[33]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_33),
        .out_chan_dep_data(out_chan_dep_data_33),
        .token_out_vec(token_out_vec_33),
        .dl_detect_out(dl_in_vec[33]));

    assign proc_33_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_27_blk_n) | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_27_blk_n) | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_WriteC_Flattened_fu_179.cPipes_27_blk_n);
    assign proc_33_data_PIPO_blk[0] = 1'b0;
    assign proc_33_start_FIFO_blk[0] = 1'b0;
    assign proc_33_TLF_FIFO_blk[0] = 1'b0;
    assign proc_33_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_33_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_33[0] = dl_detect_out ? proc_dep_vld_vec_33_reg[0] : (proc_33_data_FIFO_blk[0] | proc_33_data_PIPO_blk[0] | proc_33_start_FIFO_blk[0] | proc_33_TLF_FIFO_blk[0] | proc_33_input_sync_blk[0] | proc_33_output_sync_blk[0]);
    assign proc_33_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_28_blk_n) | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_28_blk_n) | (~ProcessingElement_28_U0.grp_ProcessingElement_28_Pipeline_WriteC_Flattened_fu_179.cPipes_28_blk_n);
    assign proc_33_data_PIPO_blk[1] = 1'b0;
    assign proc_33_start_FIFO_blk[1] = 1'b0;
    assign proc_33_TLF_FIFO_blk[1] = 1'b0;
    assign proc_33_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_33_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_33[1] = dl_detect_out ? proc_dep_vld_vec_33_reg[1] : (proc_33_data_FIFO_blk[1] | proc_33_data_PIPO_blk[1] | proc_33_start_FIFO_blk[1] | proc_33_TLF_FIFO_blk[1] | proc_33_input_sync_blk[1] | proc_33_output_sync_blk[1]);
    assign proc_33_data_FIFO_blk[2] = 1'b0;
    assign proc_33_data_PIPO_blk[2] = 1'b0;
    assign proc_33_start_FIFO_blk[2] = 1'b0;
    assign proc_33_TLF_FIFO_blk[2] = 1'b0;
    assign proc_33_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_33_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_33[2] = dl_detect_out ? proc_dep_vld_vec_33_reg[2] : (proc_33_data_FIFO_blk[2] | proc_33_data_PIPO_blk[2] | proc_33_start_FIFO_blk[2] | proc_33_TLF_FIFO_blk[2] | proc_33_input_sync_blk[2] | proc_33_output_sync_blk[2]);
    assign proc_33_data_FIFO_blk[3] = 1'b0;
    assign proc_33_data_PIPO_blk[3] = 1'b0;
    assign proc_33_start_FIFO_blk[3] = 1'b0;
    assign proc_33_TLF_FIFO_blk[3] = 1'b0;
    assign proc_33_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_33_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_33[3] = dl_detect_out ? proc_dep_vld_vec_33_reg[3] : (proc_33_data_FIFO_blk[3] | proc_33_data_PIPO_blk[3] | proc_33_start_FIFO_blk[3] | proc_33_TLF_FIFO_blk[3] | proc_33_input_sync_blk[3] | proc_33_output_sync_blk[3]);
    assign proc_33_data_FIFO_blk[4] = 1'b0;
    assign proc_33_data_PIPO_blk[4] = 1'b0;
    assign proc_33_start_FIFO_blk[4] = 1'b0;
    assign proc_33_TLF_FIFO_blk[4] = 1'b0;
    assign proc_33_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_33_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_33[4] = dl_detect_out ? proc_dep_vld_vec_33_reg[4] : (proc_33_data_FIFO_blk[4] | proc_33_data_PIPO_blk[4] | proc_33_start_FIFO_blk[4] | proc_33_TLF_FIFO_blk[4] | proc_33_input_sync_blk[4] | proc_33_output_sync_blk[4]);
    assign proc_33_data_FIFO_blk[5] = 1'b0;
    assign proc_33_data_PIPO_blk[5] = 1'b0;
    assign proc_33_start_FIFO_blk[5] = 1'b0;
    assign proc_33_TLF_FIFO_blk[5] = 1'b0;
    assign proc_33_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_33_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_33[5] = dl_detect_out ? proc_dep_vld_vec_33_reg[5] : (proc_33_data_FIFO_blk[5] | proc_33_data_PIPO_blk[5] | proc_33_start_FIFO_blk[5] | proc_33_TLF_FIFO_blk[5] | proc_33_input_sync_blk[5] | proc_33_output_sync_blk[5]);
    assign proc_33_data_FIFO_blk[6] = 1'b0;
    assign proc_33_data_PIPO_blk[6] = 1'b0;
    assign proc_33_start_FIFO_blk[6] = 1'b0;
    assign proc_33_TLF_FIFO_blk[6] = 1'b0;
    assign proc_33_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_33_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_33[6] = dl_detect_out ? proc_dep_vld_vec_33_reg[6] : (proc_33_data_FIFO_blk[6] | proc_33_data_PIPO_blk[6] | proc_33_start_FIFO_blk[6] | proc_33_TLF_FIFO_blk[6] | proc_33_input_sync_blk[6] | proc_33_output_sync_blk[6]);
    assign proc_33_data_FIFO_blk[7] = 1'b0;
    assign proc_33_data_PIPO_blk[7] = 1'b0;
    assign proc_33_start_FIFO_blk[7] = 1'b0;
    assign proc_33_TLF_FIFO_blk[7] = 1'b0;
    assign proc_33_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_33_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_33[7] = dl_detect_out ? proc_dep_vld_vec_33_reg[7] : (proc_33_data_FIFO_blk[7] | proc_33_data_PIPO_blk[7] | proc_33_start_FIFO_blk[7] | proc_33_TLF_FIFO_blk[7] | proc_33_input_sync_blk[7] | proc_33_output_sync_blk[7]);
    assign proc_33_data_FIFO_blk[8] = 1'b0;
    assign proc_33_data_PIPO_blk[8] = 1'b0;
    assign proc_33_start_FIFO_blk[8] = 1'b0;
    assign proc_33_TLF_FIFO_blk[8] = 1'b0;
    assign proc_33_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_33_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_33[8] = dl_detect_out ? proc_dep_vld_vec_33_reg[8] : (proc_33_data_FIFO_blk[8] | proc_33_data_PIPO_blk[8] | proc_33_start_FIFO_blk[8] | proc_33_TLF_FIFO_blk[8] | proc_33_input_sync_blk[8] | proc_33_output_sync_blk[8]);
    assign proc_33_data_FIFO_blk[9] = 1'b0;
    assign proc_33_data_PIPO_blk[9] = 1'b0;
    assign proc_33_start_FIFO_blk[9] = 1'b0;
    assign proc_33_TLF_FIFO_blk[9] = 1'b0;
    assign proc_33_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_33_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_33[9] = dl_detect_out ? proc_dep_vld_vec_33_reg[9] : (proc_33_data_FIFO_blk[9] | proc_33_data_PIPO_blk[9] | proc_33_start_FIFO_blk[9] | proc_33_TLF_FIFO_blk[9] | proc_33_input_sync_blk[9] | proc_33_output_sync_blk[9]);
    assign proc_33_data_FIFO_blk[10] = 1'b0;
    assign proc_33_data_PIPO_blk[10] = 1'b0;
    assign proc_33_start_FIFO_blk[10] = 1'b0;
    assign proc_33_TLF_FIFO_blk[10] = 1'b0;
    assign proc_33_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_33_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_33[10] = dl_detect_out ? proc_dep_vld_vec_33_reg[10] : (proc_33_data_FIFO_blk[10] | proc_33_data_PIPO_blk[10] | proc_33_start_FIFO_blk[10] | proc_33_TLF_FIFO_blk[10] | proc_33_input_sync_blk[10] | proc_33_output_sync_blk[10]);
    assign proc_33_data_FIFO_blk[11] = 1'b0;
    assign proc_33_data_PIPO_blk[11] = 1'b0;
    assign proc_33_start_FIFO_blk[11] = 1'b0;
    assign proc_33_TLF_FIFO_blk[11] = 1'b0;
    assign proc_33_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_33_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_33[11] = dl_detect_out ? proc_dep_vld_vec_33_reg[11] : (proc_33_data_FIFO_blk[11] | proc_33_data_PIPO_blk[11] | proc_33_start_FIFO_blk[11] | proc_33_TLF_FIFO_blk[11] | proc_33_input_sync_blk[11] | proc_33_output_sync_blk[11]);
    assign proc_33_data_FIFO_blk[12] = 1'b0;
    assign proc_33_data_PIPO_blk[12] = 1'b0;
    assign proc_33_start_FIFO_blk[12] = 1'b0;
    assign proc_33_TLF_FIFO_blk[12] = 1'b0;
    assign proc_33_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_33_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_33[12] = dl_detect_out ? proc_dep_vld_vec_33_reg[12] : (proc_33_data_FIFO_blk[12] | proc_33_data_PIPO_blk[12] | proc_33_start_FIFO_blk[12] | proc_33_TLF_FIFO_blk[12] | proc_33_input_sync_blk[12] | proc_33_output_sync_blk[12]);
    assign proc_33_data_FIFO_blk[13] = 1'b0;
    assign proc_33_data_PIPO_blk[13] = 1'b0;
    assign proc_33_start_FIFO_blk[13] = 1'b0;
    assign proc_33_TLF_FIFO_blk[13] = 1'b0;
    assign proc_33_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_33_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_33[13] = dl_detect_out ? proc_dep_vld_vec_33_reg[13] : (proc_33_data_FIFO_blk[13] | proc_33_data_PIPO_blk[13] | proc_33_start_FIFO_blk[13] | proc_33_TLF_FIFO_blk[13] | proc_33_input_sync_blk[13] | proc_33_output_sync_blk[13]);
    assign proc_33_data_FIFO_blk[14] = 1'b0;
    assign proc_33_data_PIPO_blk[14] = 1'b0;
    assign proc_33_start_FIFO_blk[14] = 1'b0;
    assign proc_33_TLF_FIFO_blk[14] = 1'b0;
    assign proc_33_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_33_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_33[14] = dl_detect_out ? proc_dep_vld_vec_33_reg[14] : (proc_33_data_FIFO_blk[14] | proc_33_data_PIPO_blk[14] | proc_33_start_FIFO_blk[14] | proc_33_TLF_FIFO_blk[14] | proc_33_input_sync_blk[14] | proc_33_output_sync_blk[14]);
    assign proc_33_data_FIFO_blk[15] = 1'b0;
    assign proc_33_data_PIPO_blk[15] = 1'b0;
    assign proc_33_start_FIFO_blk[15] = 1'b0;
    assign proc_33_TLF_FIFO_blk[15] = 1'b0;
    assign proc_33_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_33_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_33[15] = dl_detect_out ? proc_dep_vld_vec_33_reg[15] : (proc_33_data_FIFO_blk[15] | proc_33_data_PIPO_blk[15] | proc_33_start_FIFO_blk[15] | proc_33_TLF_FIFO_blk[15] | proc_33_input_sync_blk[15] | proc_33_output_sync_blk[15]);
    assign proc_33_data_FIFO_blk[16] = 1'b0;
    assign proc_33_data_PIPO_blk[16] = 1'b0;
    assign proc_33_start_FIFO_blk[16] = 1'b0;
    assign proc_33_TLF_FIFO_blk[16] = 1'b0;
    assign proc_33_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_33_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_33[16] = dl_detect_out ? proc_dep_vld_vec_33_reg[16] : (proc_33_data_FIFO_blk[16] | proc_33_data_PIPO_blk[16] | proc_33_start_FIFO_blk[16] | proc_33_TLF_FIFO_blk[16] | proc_33_input_sync_blk[16] | proc_33_output_sync_blk[16]);
    assign proc_33_data_FIFO_blk[17] = 1'b0;
    assign proc_33_data_PIPO_blk[17] = 1'b0;
    assign proc_33_start_FIFO_blk[17] = 1'b0;
    assign proc_33_TLF_FIFO_blk[17] = 1'b0;
    assign proc_33_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_33_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_33[17] = dl_detect_out ? proc_dep_vld_vec_33_reg[17] : (proc_33_data_FIFO_blk[17] | proc_33_data_PIPO_blk[17] | proc_33_start_FIFO_blk[17] | proc_33_TLF_FIFO_blk[17] | proc_33_input_sync_blk[17] | proc_33_output_sync_blk[17]);
    assign proc_33_data_FIFO_blk[18] = 1'b0;
    assign proc_33_data_PIPO_blk[18] = 1'b0;
    assign proc_33_start_FIFO_blk[18] = 1'b0;
    assign proc_33_TLF_FIFO_blk[18] = 1'b0;
    assign proc_33_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_33_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_33[18] = dl_detect_out ? proc_dep_vld_vec_33_reg[18] : (proc_33_data_FIFO_blk[18] | proc_33_data_PIPO_blk[18] | proc_33_start_FIFO_blk[18] | proc_33_TLF_FIFO_blk[18] | proc_33_input_sync_blk[18] | proc_33_output_sync_blk[18]);
    assign proc_33_data_FIFO_blk[19] = 1'b0;
    assign proc_33_data_PIPO_blk[19] = 1'b0;
    assign proc_33_start_FIFO_blk[19] = 1'b0;
    assign proc_33_TLF_FIFO_blk[19] = 1'b0;
    assign proc_33_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_33_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_33[19] = dl_detect_out ? proc_dep_vld_vec_33_reg[19] : (proc_33_data_FIFO_blk[19] | proc_33_data_PIPO_blk[19] | proc_33_start_FIFO_blk[19] | proc_33_TLF_FIFO_blk[19] | proc_33_input_sync_blk[19] | proc_33_output_sync_blk[19]);
    assign proc_33_data_FIFO_blk[20] = 1'b0;
    assign proc_33_data_PIPO_blk[20] = 1'b0;
    assign proc_33_start_FIFO_blk[20] = 1'b0;
    assign proc_33_TLF_FIFO_blk[20] = 1'b0;
    assign proc_33_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_33_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_33[20] = dl_detect_out ? proc_dep_vld_vec_33_reg[20] : (proc_33_data_FIFO_blk[20] | proc_33_data_PIPO_blk[20] | proc_33_start_FIFO_blk[20] | proc_33_TLF_FIFO_blk[20] | proc_33_input_sync_blk[20] | proc_33_output_sync_blk[20]);
    assign proc_33_data_FIFO_blk[21] = 1'b0;
    assign proc_33_data_PIPO_blk[21] = 1'b0;
    assign proc_33_start_FIFO_blk[21] = 1'b0;
    assign proc_33_TLF_FIFO_blk[21] = 1'b0;
    assign proc_33_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_33_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_33[21] = dl_detect_out ? proc_dep_vld_vec_33_reg[21] : (proc_33_data_FIFO_blk[21] | proc_33_data_PIPO_blk[21] | proc_33_start_FIFO_blk[21] | proc_33_TLF_FIFO_blk[21] | proc_33_input_sync_blk[21] | proc_33_output_sync_blk[21]);
    assign proc_33_data_FIFO_blk[22] = 1'b0;
    assign proc_33_data_PIPO_blk[22] = 1'b0;
    assign proc_33_start_FIFO_blk[22] = 1'b0;
    assign proc_33_TLF_FIFO_blk[22] = 1'b0;
    assign proc_33_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_33_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_33[22] = dl_detect_out ? proc_dep_vld_vec_33_reg[22] : (proc_33_data_FIFO_blk[22] | proc_33_data_PIPO_blk[22] | proc_33_start_FIFO_blk[22] | proc_33_TLF_FIFO_blk[22] | proc_33_input_sync_blk[22] | proc_33_output_sync_blk[22]);
    assign proc_33_data_FIFO_blk[23] = 1'b0;
    assign proc_33_data_PIPO_blk[23] = 1'b0;
    assign proc_33_start_FIFO_blk[23] = 1'b0;
    assign proc_33_TLF_FIFO_blk[23] = 1'b0;
    assign proc_33_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_33_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_33[23] = dl_detect_out ? proc_dep_vld_vec_33_reg[23] : (proc_33_data_FIFO_blk[23] | proc_33_data_PIPO_blk[23] | proc_33_start_FIFO_blk[23] | proc_33_TLF_FIFO_blk[23] | proc_33_input_sync_blk[23] | proc_33_output_sync_blk[23]);
    assign proc_33_data_FIFO_blk[24] = 1'b0;
    assign proc_33_data_PIPO_blk[24] = 1'b0;
    assign proc_33_start_FIFO_blk[24] = 1'b0;
    assign proc_33_TLF_FIFO_blk[24] = 1'b0;
    assign proc_33_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_33_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_33[24] = dl_detect_out ? proc_dep_vld_vec_33_reg[24] : (proc_33_data_FIFO_blk[24] | proc_33_data_PIPO_blk[24] | proc_33_start_FIFO_blk[24] | proc_33_TLF_FIFO_blk[24] | proc_33_input_sync_blk[24] | proc_33_output_sync_blk[24]);
    assign proc_33_data_FIFO_blk[25] = 1'b0;
    assign proc_33_data_PIPO_blk[25] = 1'b0;
    assign proc_33_start_FIFO_blk[25] = 1'b0;
    assign proc_33_TLF_FIFO_blk[25] = 1'b0;
    assign proc_33_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_33_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_33[25] = dl_detect_out ? proc_dep_vld_vec_33_reg[25] : (proc_33_data_FIFO_blk[25] | proc_33_data_PIPO_blk[25] | proc_33_start_FIFO_blk[25] | proc_33_TLF_FIFO_blk[25] | proc_33_input_sync_blk[25] | proc_33_output_sync_blk[25]);
    assign proc_33_data_FIFO_blk[26] = 1'b0;
    assign proc_33_data_PIPO_blk[26] = 1'b0;
    assign proc_33_start_FIFO_blk[26] = 1'b0;
    assign proc_33_TLF_FIFO_blk[26] = 1'b0;
    assign proc_33_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_33_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_33[26] = dl_detect_out ? proc_dep_vld_vec_33_reg[26] : (proc_33_data_FIFO_blk[26] | proc_33_data_PIPO_blk[26] | proc_33_start_FIFO_blk[26] | proc_33_TLF_FIFO_blk[26] | proc_33_input_sync_blk[26] | proc_33_output_sync_blk[26]);
    assign proc_33_data_FIFO_blk[27] = 1'b0;
    assign proc_33_data_PIPO_blk[27] = 1'b0;
    assign proc_33_start_FIFO_blk[27] = 1'b0;
    assign proc_33_TLF_FIFO_blk[27] = 1'b0;
    assign proc_33_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_33_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_33[27] = dl_detect_out ? proc_dep_vld_vec_33_reg[27] : (proc_33_data_FIFO_blk[27] | proc_33_data_PIPO_blk[27] | proc_33_start_FIFO_blk[27] | proc_33_TLF_FIFO_blk[27] | proc_33_input_sync_blk[27] | proc_33_output_sync_blk[27]);
    assign proc_33_data_FIFO_blk[28] = 1'b0;
    assign proc_33_data_PIPO_blk[28] = 1'b0;
    assign proc_33_start_FIFO_blk[28] = 1'b0;
    assign proc_33_TLF_FIFO_blk[28] = 1'b0;
    assign proc_33_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_33_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_33[28] = dl_detect_out ? proc_dep_vld_vec_33_reg[28] : (proc_33_data_FIFO_blk[28] | proc_33_data_PIPO_blk[28] | proc_33_start_FIFO_blk[28] | proc_33_TLF_FIFO_blk[28] | proc_33_input_sync_blk[28] | proc_33_output_sync_blk[28]);
    assign proc_33_data_FIFO_blk[29] = 1'b0;
    assign proc_33_data_PIPO_blk[29] = 1'b0;
    assign proc_33_start_FIFO_blk[29] = 1'b0;
    assign proc_33_TLF_FIFO_blk[29] = 1'b0;
    assign proc_33_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_33_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_33[29] = dl_detect_out ? proc_dep_vld_vec_33_reg[29] : (proc_33_data_FIFO_blk[29] | proc_33_data_PIPO_blk[29] | proc_33_start_FIFO_blk[29] | proc_33_TLF_FIFO_blk[29] | proc_33_input_sync_blk[29] | proc_33_output_sync_blk[29]);
    assign proc_33_data_FIFO_blk[30] = 1'b0;
    assign proc_33_data_PIPO_blk[30] = 1'b0;
    assign proc_33_start_FIFO_blk[30] = 1'b0;
    assign proc_33_TLF_FIFO_blk[30] = 1'b0;
    assign proc_33_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_33_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_33[30] = dl_detect_out ? proc_dep_vld_vec_33_reg[30] : (proc_33_data_FIFO_blk[30] | proc_33_data_PIPO_blk[30] | proc_33_start_FIFO_blk[30] | proc_33_TLF_FIFO_blk[30] | proc_33_input_sync_blk[30] | proc_33_output_sync_blk[30]);
    assign proc_33_data_FIFO_blk[31] = 1'b0;
    assign proc_33_data_PIPO_blk[31] = 1'b0;
    assign proc_33_start_FIFO_blk[31] = 1'b0;
    assign proc_33_TLF_FIFO_blk[31] = 1'b0;
    assign proc_33_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_33_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_33[31] = dl_detect_out ? proc_dep_vld_vec_33_reg[31] : (proc_33_data_FIFO_blk[31] | proc_33_data_PIPO_blk[31] | proc_33_start_FIFO_blk[31] | proc_33_TLF_FIFO_blk[31] | proc_33_input_sync_blk[31] | proc_33_output_sync_blk[31]);
    assign proc_33_data_FIFO_blk[32] = 1'b0;
    assign proc_33_data_PIPO_blk[32] = 1'b0;
    assign proc_33_start_FIFO_blk[32] = 1'b0;
    assign proc_33_TLF_FIFO_blk[32] = 1'b0;
    assign proc_33_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_28_U0_ap_ready & ProcessingElement_28_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_33_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_33[32] = dl_detect_out ? proc_dep_vld_vec_33_reg[32] : (proc_33_data_FIFO_blk[32] | proc_33_data_PIPO_blk[32] | proc_33_start_FIFO_blk[32] | proc_33_TLF_FIFO_blk[32] | proc_33_input_sync_blk[32] | proc_33_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_33_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_33_reg <= proc_dep_vld_vec_33;
        end
    end
    assign in_chan_dep_vld_vec_33[0] = dep_chan_vld_0_33;
    assign in_chan_dep_data_vec_33[39 : 0] = dep_chan_data_0_33;
    assign token_in_vec_33[0] = token_0_33;
    assign in_chan_dep_vld_vec_33[1] = dep_chan_vld_1_33;
    assign in_chan_dep_data_vec_33[79 : 40] = dep_chan_data_1_33;
    assign token_in_vec_33[1] = token_1_33;
    assign in_chan_dep_vld_vec_33[2] = dep_chan_vld_3_33;
    assign in_chan_dep_data_vec_33[119 : 80] = dep_chan_data_3_33;
    assign token_in_vec_33[2] = token_3_33;
    assign in_chan_dep_vld_vec_33[3] = dep_chan_vld_6_33;
    assign in_chan_dep_data_vec_33[159 : 120] = dep_chan_data_6_33;
    assign token_in_vec_33[3] = token_6_33;
    assign in_chan_dep_vld_vec_33[4] = dep_chan_vld_7_33;
    assign in_chan_dep_data_vec_33[199 : 160] = dep_chan_data_7_33;
    assign token_in_vec_33[4] = token_7_33;
    assign in_chan_dep_vld_vec_33[5] = dep_chan_vld_8_33;
    assign in_chan_dep_data_vec_33[239 : 200] = dep_chan_data_8_33;
    assign token_in_vec_33[5] = token_8_33;
    assign in_chan_dep_vld_vec_33[6] = dep_chan_vld_9_33;
    assign in_chan_dep_data_vec_33[279 : 240] = dep_chan_data_9_33;
    assign token_in_vec_33[6] = token_9_33;
    assign in_chan_dep_vld_vec_33[7] = dep_chan_vld_10_33;
    assign in_chan_dep_data_vec_33[319 : 280] = dep_chan_data_10_33;
    assign token_in_vec_33[7] = token_10_33;
    assign in_chan_dep_vld_vec_33[8] = dep_chan_vld_11_33;
    assign in_chan_dep_data_vec_33[359 : 320] = dep_chan_data_11_33;
    assign token_in_vec_33[8] = token_11_33;
    assign in_chan_dep_vld_vec_33[9] = dep_chan_vld_12_33;
    assign in_chan_dep_data_vec_33[399 : 360] = dep_chan_data_12_33;
    assign token_in_vec_33[9] = token_12_33;
    assign in_chan_dep_vld_vec_33[10] = dep_chan_vld_13_33;
    assign in_chan_dep_data_vec_33[439 : 400] = dep_chan_data_13_33;
    assign token_in_vec_33[10] = token_13_33;
    assign in_chan_dep_vld_vec_33[11] = dep_chan_vld_14_33;
    assign in_chan_dep_data_vec_33[479 : 440] = dep_chan_data_14_33;
    assign token_in_vec_33[11] = token_14_33;
    assign in_chan_dep_vld_vec_33[12] = dep_chan_vld_15_33;
    assign in_chan_dep_data_vec_33[519 : 480] = dep_chan_data_15_33;
    assign token_in_vec_33[12] = token_15_33;
    assign in_chan_dep_vld_vec_33[13] = dep_chan_vld_16_33;
    assign in_chan_dep_data_vec_33[559 : 520] = dep_chan_data_16_33;
    assign token_in_vec_33[13] = token_16_33;
    assign in_chan_dep_vld_vec_33[14] = dep_chan_vld_17_33;
    assign in_chan_dep_data_vec_33[599 : 560] = dep_chan_data_17_33;
    assign token_in_vec_33[14] = token_17_33;
    assign in_chan_dep_vld_vec_33[15] = dep_chan_vld_18_33;
    assign in_chan_dep_data_vec_33[639 : 600] = dep_chan_data_18_33;
    assign token_in_vec_33[15] = token_18_33;
    assign in_chan_dep_vld_vec_33[16] = dep_chan_vld_19_33;
    assign in_chan_dep_data_vec_33[679 : 640] = dep_chan_data_19_33;
    assign token_in_vec_33[16] = token_19_33;
    assign in_chan_dep_vld_vec_33[17] = dep_chan_vld_20_33;
    assign in_chan_dep_data_vec_33[719 : 680] = dep_chan_data_20_33;
    assign token_in_vec_33[17] = token_20_33;
    assign in_chan_dep_vld_vec_33[18] = dep_chan_vld_21_33;
    assign in_chan_dep_data_vec_33[759 : 720] = dep_chan_data_21_33;
    assign token_in_vec_33[18] = token_21_33;
    assign in_chan_dep_vld_vec_33[19] = dep_chan_vld_22_33;
    assign in_chan_dep_data_vec_33[799 : 760] = dep_chan_data_22_33;
    assign token_in_vec_33[19] = token_22_33;
    assign in_chan_dep_vld_vec_33[20] = dep_chan_vld_23_33;
    assign in_chan_dep_data_vec_33[839 : 800] = dep_chan_data_23_33;
    assign token_in_vec_33[20] = token_23_33;
    assign in_chan_dep_vld_vec_33[21] = dep_chan_vld_24_33;
    assign in_chan_dep_data_vec_33[879 : 840] = dep_chan_data_24_33;
    assign token_in_vec_33[21] = token_24_33;
    assign in_chan_dep_vld_vec_33[22] = dep_chan_vld_25_33;
    assign in_chan_dep_data_vec_33[919 : 880] = dep_chan_data_25_33;
    assign token_in_vec_33[22] = token_25_33;
    assign in_chan_dep_vld_vec_33[23] = dep_chan_vld_26_33;
    assign in_chan_dep_data_vec_33[959 : 920] = dep_chan_data_26_33;
    assign token_in_vec_33[23] = token_26_33;
    assign in_chan_dep_vld_vec_33[24] = dep_chan_vld_27_33;
    assign in_chan_dep_data_vec_33[999 : 960] = dep_chan_data_27_33;
    assign token_in_vec_33[24] = token_27_33;
    assign in_chan_dep_vld_vec_33[25] = dep_chan_vld_28_33;
    assign in_chan_dep_data_vec_33[1039 : 1000] = dep_chan_data_28_33;
    assign token_in_vec_33[25] = token_28_33;
    assign in_chan_dep_vld_vec_33[26] = dep_chan_vld_29_33;
    assign in_chan_dep_data_vec_33[1079 : 1040] = dep_chan_data_29_33;
    assign token_in_vec_33[26] = token_29_33;
    assign in_chan_dep_vld_vec_33[27] = dep_chan_vld_30_33;
    assign in_chan_dep_data_vec_33[1119 : 1080] = dep_chan_data_30_33;
    assign token_in_vec_33[27] = token_30_33;
    assign in_chan_dep_vld_vec_33[28] = dep_chan_vld_31_33;
    assign in_chan_dep_data_vec_33[1159 : 1120] = dep_chan_data_31_33;
    assign token_in_vec_33[28] = token_31_33;
    assign in_chan_dep_vld_vec_33[29] = dep_chan_vld_32_33;
    assign in_chan_dep_data_vec_33[1199 : 1160] = dep_chan_data_32_33;
    assign token_in_vec_33[29] = token_32_33;
    assign in_chan_dep_vld_vec_33[30] = dep_chan_vld_34_33;
    assign in_chan_dep_data_vec_33[1239 : 1200] = dep_chan_data_34_33;
    assign token_in_vec_33[30] = token_34_33;
    assign in_chan_dep_vld_vec_33[31] = dep_chan_vld_35_33;
    assign in_chan_dep_data_vec_33[1279 : 1240] = dep_chan_data_35_33;
    assign token_in_vec_33[31] = token_35_33;
    assign in_chan_dep_vld_vec_33[32] = dep_chan_vld_36_33;
    assign in_chan_dep_data_vec_33[1319 : 1280] = dep_chan_data_36_33;
    assign token_in_vec_33[32] = token_36_33;
    assign dep_chan_vld_33_32 = out_chan_dep_vld_vec_33[0];
    assign dep_chan_data_33_32 = out_chan_dep_data_33;
    assign token_33_32 = token_out_vec_33[0];
    assign dep_chan_vld_33_34 = out_chan_dep_vld_vec_33[1];
    assign dep_chan_data_33_34 = out_chan_dep_data_33;
    assign token_33_34 = token_out_vec_33[1];
    assign dep_chan_vld_33_0 = out_chan_dep_vld_vec_33[2];
    assign dep_chan_data_33_0 = out_chan_dep_data_33;
    assign token_33_0 = token_out_vec_33[2];
    assign dep_chan_vld_33_1 = out_chan_dep_vld_vec_33[3];
    assign dep_chan_data_33_1 = out_chan_dep_data_33;
    assign token_33_1 = token_out_vec_33[3];
    assign dep_chan_vld_33_3 = out_chan_dep_vld_vec_33[4];
    assign dep_chan_data_33_3 = out_chan_dep_data_33;
    assign token_33_3 = token_out_vec_33[4];
    assign dep_chan_vld_33_6 = out_chan_dep_vld_vec_33[5];
    assign dep_chan_data_33_6 = out_chan_dep_data_33;
    assign token_33_6 = token_out_vec_33[5];
    assign dep_chan_vld_33_7 = out_chan_dep_vld_vec_33[6];
    assign dep_chan_data_33_7 = out_chan_dep_data_33;
    assign token_33_7 = token_out_vec_33[6];
    assign dep_chan_vld_33_8 = out_chan_dep_vld_vec_33[7];
    assign dep_chan_data_33_8 = out_chan_dep_data_33;
    assign token_33_8 = token_out_vec_33[7];
    assign dep_chan_vld_33_9 = out_chan_dep_vld_vec_33[8];
    assign dep_chan_data_33_9 = out_chan_dep_data_33;
    assign token_33_9 = token_out_vec_33[8];
    assign dep_chan_vld_33_10 = out_chan_dep_vld_vec_33[9];
    assign dep_chan_data_33_10 = out_chan_dep_data_33;
    assign token_33_10 = token_out_vec_33[9];
    assign dep_chan_vld_33_11 = out_chan_dep_vld_vec_33[10];
    assign dep_chan_data_33_11 = out_chan_dep_data_33;
    assign token_33_11 = token_out_vec_33[10];
    assign dep_chan_vld_33_12 = out_chan_dep_vld_vec_33[11];
    assign dep_chan_data_33_12 = out_chan_dep_data_33;
    assign token_33_12 = token_out_vec_33[11];
    assign dep_chan_vld_33_13 = out_chan_dep_vld_vec_33[12];
    assign dep_chan_data_33_13 = out_chan_dep_data_33;
    assign token_33_13 = token_out_vec_33[12];
    assign dep_chan_vld_33_14 = out_chan_dep_vld_vec_33[13];
    assign dep_chan_data_33_14 = out_chan_dep_data_33;
    assign token_33_14 = token_out_vec_33[13];
    assign dep_chan_vld_33_15 = out_chan_dep_vld_vec_33[14];
    assign dep_chan_data_33_15 = out_chan_dep_data_33;
    assign token_33_15 = token_out_vec_33[14];
    assign dep_chan_vld_33_16 = out_chan_dep_vld_vec_33[15];
    assign dep_chan_data_33_16 = out_chan_dep_data_33;
    assign token_33_16 = token_out_vec_33[15];
    assign dep_chan_vld_33_17 = out_chan_dep_vld_vec_33[16];
    assign dep_chan_data_33_17 = out_chan_dep_data_33;
    assign token_33_17 = token_out_vec_33[16];
    assign dep_chan_vld_33_18 = out_chan_dep_vld_vec_33[17];
    assign dep_chan_data_33_18 = out_chan_dep_data_33;
    assign token_33_18 = token_out_vec_33[17];
    assign dep_chan_vld_33_19 = out_chan_dep_vld_vec_33[18];
    assign dep_chan_data_33_19 = out_chan_dep_data_33;
    assign token_33_19 = token_out_vec_33[18];
    assign dep_chan_vld_33_20 = out_chan_dep_vld_vec_33[19];
    assign dep_chan_data_33_20 = out_chan_dep_data_33;
    assign token_33_20 = token_out_vec_33[19];
    assign dep_chan_vld_33_21 = out_chan_dep_vld_vec_33[20];
    assign dep_chan_data_33_21 = out_chan_dep_data_33;
    assign token_33_21 = token_out_vec_33[20];
    assign dep_chan_vld_33_22 = out_chan_dep_vld_vec_33[21];
    assign dep_chan_data_33_22 = out_chan_dep_data_33;
    assign token_33_22 = token_out_vec_33[21];
    assign dep_chan_vld_33_23 = out_chan_dep_vld_vec_33[22];
    assign dep_chan_data_33_23 = out_chan_dep_data_33;
    assign token_33_23 = token_out_vec_33[22];
    assign dep_chan_vld_33_24 = out_chan_dep_vld_vec_33[23];
    assign dep_chan_data_33_24 = out_chan_dep_data_33;
    assign token_33_24 = token_out_vec_33[23];
    assign dep_chan_vld_33_25 = out_chan_dep_vld_vec_33[24];
    assign dep_chan_data_33_25 = out_chan_dep_data_33;
    assign token_33_25 = token_out_vec_33[24];
    assign dep_chan_vld_33_26 = out_chan_dep_vld_vec_33[25];
    assign dep_chan_data_33_26 = out_chan_dep_data_33;
    assign token_33_26 = token_out_vec_33[25];
    assign dep_chan_vld_33_27 = out_chan_dep_vld_vec_33[26];
    assign dep_chan_data_33_27 = out_chan_dep_data_33;
    assign token_33_27 = token_out_vec_33[26];
    assign dep_chan_vld_33_28 = out_chan_dep_vld_vec_33[27];
    assign dep_chan_data_33_28 = out_chan_dep_data_33;
    assign token_33_28 = token_out_vec_33[27];
    assign dep_chan_vld_33_29 = out_chan_dep_vld_vec_33[28];
    assign dep_chan_data_33_29 = out_chan_dep_data_33;
    assign token_33_29 = token_out_vec_33[28];
    assign dep_chan_vld_33_30 = out_chan_dep_vld_vec_33[29];
    assign dep_chan_data_33_30 = out_chan_dep_data_33;
    assign token_33_30 = token_out_vec_33[29];
    assign dep_chan_vld_33_31 = out_chan_dep_vld_vec_33[30];
    assign dep_chan_data_33_31 = out_chan_dep_data_33;
    assign token_33_31 = token_out_vec_33[30];
    assign dep_chan_vld_33_35 = out_chan_dep_vld_vec_33[31];
    assign dep_chan_data_33_35 = out_chan_dep_data_33;
    assign token_33_35 = token_out_vec_33[31];
    assign dep_chan_vld_33_36 = out_chan_dep_vld_vec_33[32];
    assign dep_chan_data_33_36 = out_chan_dep_data_33;
    assign token_33_36 = token_out_vec_33[32];

    // Process: ProcessingElement_29_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 34, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_34 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_34),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_34),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_34),
        .token_in_vec(token_in_vec_34),
        .dl_detect_in(dl_detect_out),
        .origin(origin[34]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_34),
        .out_chan_dep_data(out_chan_dep_data_34),
        .token_out_vec(token_out_vec_34),
        .dl_detect_out(dl_in_vec[34]));

    assign proc_34_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_28_blk_n) | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_28_blk_n) | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_WriteC_Flattened_fu_179.cPipes_28_blk_n);
    assign proc_34_data_PIPO_blk[0] = 1'b0;
    assign proc_34_start_FIFO_blk[0] = 1'b0;
    assign proc_34_TLF_FIFO_blk[0] = 1'b0;
    assign proc_34_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_34_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_34[0] = dl_detect_out ? proc_dep_vld_vec_34_reg[0] : (proc_34_data_FIFO_blk[0] | proc_34_data_PIPO_blk[0] | proc_34_start_FIFO_blk[0] | proc_34_TLF_FIFO_blk[0] | proc_34_input_sync_blk[0] | proc_34_output_sync_blk[0]);
    assign proc_34_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_148.aPipes_29_blk_n) | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_29_blk_n) | (~ProcessingElement_29_U0.grp_ProcessingElement_29_Pipeline_WriteC_Flattened_fu_179.cPipes_29_blk_n);
    assign proc_34_data_PIPO_blk[1] = 1'b0;
    assign proc_34_start_FIFO_blk[1] = 1'b0;
    assign proc_34_TLF_FIFO_blk[1] = 1'b0;
    assign proc_34_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_34_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_34[1] = dl_detect_out ? proc_dep_vld_vec_34_reg[1] : (proc_34_data_FIFO_blk[1] | proc_34_data_PIPO_blk[1] | proc_34_start_FIFO_blk[1] | proc_34_TLF_FIFO_blk[1] | proc_34_input_sync_blk[1] | proc_34_output_sync_blk[1]);
    assign proc_34_data_FIFO_blk[2] = 1'b0;
    assign proc_34_data_PIPO_blk[2] = 1'b0;
    assign proc_34_start_FIFO_blk[2] = 1'b0;
    assign proc_34_TLF_FIFO_blk[2] = 1'b0;
    assign proc_34_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_34_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_34[2] = dl_detect_out ? proc_dep_vld_vec_34_reg[2] : (proc_34_data_FIFO_blk[2] | proc_34_data_PIPO_blk[2] | proc_34_start_FIFO_blk[2] | proc_34_TLF_FIFO_blk[2] | proc_34_input_sync_blk[2] | proc_34_output_sync_blk[2]);
    assign proc_34_data_FIFO_blk[3] = 1'b0;
    assign proc_34_data_PIPO_blk[3] = 1'b0;
    assign proc_34_start_FIFO_blk[3] = 1'b0;
    assign proc_34_TLF_FIFO_blk[3] = 1'b0;
    assign proc_34_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_34_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_34[3] = dl_detect_out ? proc_dep_vld_vec_34_reg[3] : (proc_34_data_FIFO_blk[3] | proc_34_data_PIPO_blk[3] | proc_34_start_FIFO_blk[3] | proc_34_TLF_FIFO_blk[3] | proc_34_input_sync_blk[3] | proc_34_output_sync_blk[3]);
    assign proc_34_data_FIFO_blk[4] = 1'b0;
    assign proc_34_data_PIPO_blk[4] = 1'b0;
    assign proc_34_start_FIFO_blk[4] = 1'b0;
    assign proc_34_TLF_FIFO_blk[4] = 1'b0;
    assign proc_34_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_34_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_34[4] = dl_detect_out ? proc_dep_vld_vec_34_reg[4] : (proc_34_data_FIFO_blk[4] | proc_34_data_PIPO_blk[4] | proc_34_start_FIFO_blk[4] | proc_34_TLF_FIFO_blk[4] | proc_34_input_sync_blk[4] | proc_34_output_sync_blk[4]);
    assign proc_34_data_FIFO_blk[5] = 1'b0;
    assign proc_34_data_PIPO_blk[5] = 1'b0;
    assign proc_34_start_FIFO_blk[5] = 1'b0;
    assign proc_34_TLF_FIFO_blk[5] = 1'b0;
    assign proc_34_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_34_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_34[5] = dl_detect_out ? proc_dep_vld_vec_34_reg[5] : (proc_34_data_FIFO_blk[5] | proc_34_data_PIPO_blk[5] | proc_34_start_FIFO_blk[5] | proc_34_TLF_FIFO_blk[5] | proc_34_input_sync_blk[5] | proc_34_output_sync_blk[5]);
    assign proc_34_data_FIFO_blk[6] = 1'b0;
    assign proc_34_data_PIPO_blk[6] = 1'b0;
    assign proc_34_start_FIFO_blk[6] = 1'b0;
    assign proc_34_TLF_FIFO_blk[6] = 1'b0;
    assign proc_34_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_34_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_34[6] = dl_detect_out ? proc_dep_vld_vec_34_reg[6] : (proc_34_data_FIFO_blk[6] | proc_34_data_PIPO_blk[6] | proc_34_start_FIFO_blk[6] | proc_34_TLF_FIFO_blk[6] | proc_34_input_sync_blk[6] | proc_34_output_sync_blk[6]);
    assign proc_34_data_FIFO_blk[7] = 1'b0;
    assign proc_34_data_PIPO_blk[7] = 1'b0;
    assign proc_34_start_FIFO_blk[7] = 1'b0;
    assign proc_34_TLF_FIFO_blk[7] = 1'b0;
    assign proc_34_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_34_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_34[7] = dl_detect_out ? proc_dep_vld_vec_34_reg[7] : (proc_34_data_FIFO_blk[7] | proc_34_data_PIPO_blk[7] | proc_34_start_FIFO_blk[7] | proc_34_TLF_FIFO_blk[7] | proc_34_input_sync_blk[7] | proc_34_output_sync_blk[7]);
    assign proc_34_data_FIFO_blk[8] = 1'b0;
    assign proc_34_data_PIPO_blk[8] = 1'b0;
    assign proc_34_start_FIFO_blk[8] = 1'b0;
    assign proc_34_TLF_FIFO_blk[8] = 1'b0;
    assign proc_34_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_34_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_34[8] = dl_detect_out ? proc_dep_vld_vec_34_reg[8] : (proc_34_data_FIFO_blk[8] | proc_34_data_PIPO_blk[8] | proc_34_start_FIFO_blk[8] | proc_34_TLF_FIFO_blk[8] | proc_34_input_sync_blk[8] | proc_34_output_sync_blk[8]);
    assign proc_34_data_FIFO_blk[9] = 1'b0;
    assign proc_34_data_PIPO_blk[9] = 1'b0;
    assign proc_34_start_FIFO_blk[9] = 1'b0;
    assign proc_34_TLF_FIFO_blk[9] = 1'b0;
    assign proc_34_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_34_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_34[9] = dl_detect_out ? proc_dep_vld_vec_34_reg[9] : (proc_34_data_FIFO_blk[9] | proc_34_data_PIPO_blk[9] | proc_34_start_FIFO_blk[9] | proc_34_TLF_FIFO_blk[9] | proc_34_input_sync_blk[9] | proc_34_output_sync_blk[9]);
    assign proc_34_data_FIFO_blk[10] = 1'b0;
    assign proc_34_data_PIPO_blk[10] = 1'b0;
    assign proc_34_start_FIFO_blk[10] = 1'b0;
    assign proc_34_TLF_FIFO_blk[10] = 1'b0;
    assign proc_34_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_34_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_34[10] = dl_detect_out ? proc_dep_vld_vec_34_reg[10] : (proc_34_data_FIFO_blk[10] | proc_34_data_PIPO_blk[10] | proc_34_start_FIFO_blk[10] | proc_34_TLF_FIFO_blk[10] | proc_34_input_sync_blk[10] | proc_34_output_sync_blk[10]);
    assign proc_34_data_FIFO_blk[11] = 1'b0;
    assign proc_34_data_PIPO_blk[11] = 1'b0;
    assign proc_34_start_FIFO_blk[11] = 1'b0;
    assign proc_34_TLF_FIFO_blk[11] = 1'b0;
    assign proc_34_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_34_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_34[11] = dl_detect_out ? proc_dep_vld_vec_34_reg[11] : (proc_34_data_FIFO_blk[11] | proc_34_data_PIPO_blk[11] | proc_34_start_FIFO_blk[11] | proc_34_TLF_FIFO_blk[11] | proc_34_input_sync_blk[11] | proc_34_output_sync_blk[11]);
    assign proc_34_data_FIFO_blk[12] = 1'b0;
    assign proc_34_data_PIPO_blk[12] = 1'b0;
    assign proc_34_start_FIFO_blk[12] = 1'b0;
    assign proc_34_TLF_FIFO_blk[12] = 1'b0;
    assign proc_34_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_34_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_34[12] = dl_detect_out ? proc_dep_vld_vec_34_reg[12] : (proc_34_data_FIFO_blk[12] | proc_34_data_PIPO_blk[12] | proc_34_start_FIFO_blk[12] | proc_34_TLF_FIFO_blk[12] | proc_34_input_sync_blk[12] | proc_34_output_sync_blk[12]);
    assign proc_34_data_FIFO_blk[13] = 1'b0;
    assign proc_34_data_PIPO_blk[13] = 1'b0;
    assign proc_34_start_FIFO_blk[13] = 1'b0;
    assign proc_34_TLF_FIFO_blk[13] = 1'b0;
    assign proc_34_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_34_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_34[13] = dl_detect_out ? proc_dep_vld_vec_34_reg[13] : (proc_34_data_FIFO_blk[13] | proc_34_data_PIPO_blk[13] | proc_34_start_FIFO_blk[13] | proc_34_TLF_FIFO_blk[13] | proc_34_input_sync_blk[13] | proc_34_output_sync_blk[13]);
    assign proc_34_data_FIFO_blk[14] = 1'b0;
    assign proc_34_data_PIPO_blk[14] = 1'b0;
    assign proc_34_start_FIFO_blk[14] = 1'b0;
    assign proc_34_TLF_FIFO_blk[14] = 1'b0;
    assign proc_34_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_34_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_34[14] = dl_detect_out ? proc_dep_vld_vec_34_reg[14] : (proc_34_data_FIFO_blk[14] | proc_34_data_PIPO_blk[14] | proc_34_start_FIFO_blk[14] | proc_34_TLF_FIFO_blk[14] | proc_34_input_sync_blk[14] | proc_34_output_sync_blk[14]);
    assign proc_34_data_FIFO_blk[15] = 1'b0;
    assign proc_34_data_PIPO_blk[15] = 1'b0;
    assign proc_34_start_FIFO_blk[15] = 1'b0;
    assign proc_34_TLF_FIFO_blk[15] = 1'b0;
    assign proc_34_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_34_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_34[15] = dl_detect_out ? proc_dep_vld_vec_34_reg[15] : (proc_34_data_FIFO_blk[15] | proc_34_data_PIPO_blk[15] | proc_34_start_FIFO_blk[15] | proc_34_TLF_FIFO_blk[15] | proc_34_input_sync_blk[15] | proc_34_output_sync_blk[15]);
    assign proc_34_data_FIFO_blk[16] = 1'b0;
    assign proc_34_data_PIPO_blk[16] = 1'b0;
    assign proc_34_start_FIFO_blk[16] = 1'b0;
    assign proc_34_TLF_FIFO_blk[16] = 1'b0;
    assign proc_34_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_34_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_34[16] = dl_detect_out ? proc_dep_vld_vec_34_reg[16] : (proc_34_data_FIFO_blk[16] | proc_34_data_PIPO_blk[16] | proc_34_start_FIFO_blk[16] | proc_34_TLF_FIFO_blk[16] | proc_34_input_sync_blk[16] | proc_34_output_sync_blk[16]);
    assign proc_34_data_FIFO_blk[17] = 1'b0;
    assign proc_34_data_PIPO_blk[17] = 1'b0;
    assign proc_34_start_FIFO_blk[17] = 1'b0;
    assign proc_34_TLF_FIFO_blk[17] = 1'b0;
    assign proc_34_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_34_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_34[17] = dl_detect_out ? proc_dep_vld_vec_34_reg[17] : (proc_34_data_FIFO_blk[17] | proc_34_data_PIPO_blk[17] | proc_34_start_FIFO_blk[17] | proc_34_TLF_FIFO_blk[17] | proc_34_input_sync_blk[17] | proc_34_output_sync_blk[17]);
    assign proc_34_data_FIFO_blk[18] = 1'b0;
    assign proc_34_data_PIPO_blk[18] = 1'b0;
    assign proc_34_start_FIFO_blk[18] = 1'b0;
    assign proc_34_TLF_FIFO_blk[18] = 1'b0;
    assign proc_34_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_34_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_34[18] = dl_detect_out ? proc_dep_vld_vec_34_reg[18] : (proc_34_data_FIFO_blk[18] | proc_34_data_PIPO_blk[18] | proc_34_start_FIFO_blk[18] | proc_34_TLF_FIFO_blk[18] | proc_34_input_sync_blk[18] | proc_34_output_sync_blk[18]);
    assign proc_34_data_FIFO_blk[19] = 1'b0;
    assign proc_34_data_PIPO_blk[19] = 1'b0;
    assign proc_34_start_FIFO_blk[19] = 1'b0;
    assign proc_34_TLF_FIFO_blk[19] = 1'b0;
    assign proc_34_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_34_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_34[19] = dl_detect_out ? proc_dep_vld_vec_34_reg[19] : (proc_34_data_FIFO_blk[19] | proc_34_data_PIPO_blk[19] | proc_34_start_FIFO_blk[19] | proc_34_TLF_FIFO_blk[19] | proc_34_input_sync_blk[19] | proc_34_output_sync_blk[19]);
    assign proc_34_data_FIFO_blk[20] = 1'b0;
    assign proc_34_data_PIPO_blk[20] = 1'b0;
    assign proc_34_start_FIFO_blk[20] = 1'b0;
    assign proc_34_TLF_FIFO_blk[20] = 1'b0;
    assign proc_34_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_34_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_34[20] = dl_detect_out ? proc_dep_vld_vec_34_reg[20] : (proc_34_data_FIFO_blk[20] | proc_34_data_PIPO_blk[20] | proc_34_start_FIFO_blk[20] | proc_34_TLF_FIFO_blk[20] | proc_34_input_sync_blk[20] | proc_34_output_sync_blk[20]);
    assign proc_34_data_FIFO_blk[21] = 1'b0;
    assign proc_34_data_PIPO_blk[21] = 1'b0;
    assign proc_34_start_FIFO_blk[21] = 1'b0;
    assign proc_34_TLF_FIFO_blk[21] = 1'b0;
    assign proc_34_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_34_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_34[21] = dl_detect_out ? proc_dep_vld_vec_34_reg[21] : (proc_34_data_FIFO_blk[21] | proc_34_data_PIPO_blk[21] | proc_34_start_FIFO_blk[21] | proc_34_TLF_FIFO_blk[21] | proc_34_input_sync_blk[21] | proc_34_output_sync_blk[21]);
    assign proc_34_data_FIFO_blk[22] = 1'b0;
    assign proc_34_data_PIPO_blk[22] = 1'b0;
    assign proc_34_start_FIFO_blk[22] = 1'b0;
    assign proc_34_TLF_FIFO_blk[22] = 1'b0;
    assign proc_34_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_34_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_34[22] = dl_detect_out ? proc_dep_vld_vec_34_reg[22] : (proc_34_data_FIFO_blk[22] | proc_34_data_PIPO_blk[22] | proc_34_start_FIFO_blk[22] | proc_34_TLF_FIFO_blk[22] | proc_34_input_sync_blk[22] | proc_34_output_sync_blk[22]);
    assign proc_34_data_FIFO_blk[23] = 1'b0;
    assign proc_34_data_PIPO_blk[23] = 1'b0;
    assign proc_34_start_FIFO_blk[23] = 1'b0;
    assign proc_34_TLF_FIFO_blk[23] = 1'b0;
    assign proc_34_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_34_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_34[23] = dl_detect_out ? proc_dep_vld_vec_34_reg[23] : (proc_34_data_FIFO_blk[23] | proc_34_data_PIPO_blk[23] | proc_34_start_FIFO_blk[23] | proc_34_TLF_FIFO_blk[23] | proc_34_input_sync_blk[23] | proc_34_output_sync_blk[23]);
    assign proc_34_data_FIFO_blk[24] = 1'b0;
    assign proc_34_data_PIPO_blk[24] = 1'b0;
    assign proc_34_start_FIFO_blk[24] = 1'b0;
    assign proc_34_TLF_FIFO_blk[24] = 1'b0;
    assign proc_34_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_34_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_34[24] = dl_detect_out ? proc_dep_vld_vec_34_reg[24] : (proc_34_data_FIFO_blk[24] | proc_34_data_PIPO_blk[24] | proc_34_start_FIFO_blk[24] | proc_34_TLF_FIFO_blk[24] | proc_34_input_sync_blk[24] | proc_34_output_sync_blk[24]);
    assign proc_34_data_FIFO_blk[25] = 1'b0;
    assign proc_34_data_PIPO_blk[25] = 1'b0;
    assign proc_34_start_FIFO_blk[25] = 1'b0;
    assign proc_34_TLF_FIFO_blk[25] = 1'b0;
    assign proc_34_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_34_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_34[25] = dl_detect_out ? proc_dep_vld_vec_34_reg[25] : (proc_34_data_FIFO_blk[25] | proc_34_data_PIPO_blk[25] | proc_34_start_FIFO_blk[25] | proc_34_TLF_FIFO_blk[25] | proc_34_input_sync_blk[25] | proc_34_output_sync_blk[25]);
    assign proc_34_data_FIFO_blk[26] = 1'b0;
    assign proc_34_data_PIPO_blk[26] = 1'b0;
    assign proc_34_start_FIFO_blk[26] = 1'b0;
    assign proc_34_TLF_FIFO_blk[26] = 1'b0;
    assign proc_34_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_34_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_34[26] = dl_detect_out ? proc_dep_vld_vec_34_reg[26] : (proc_34_data_FIFO_blk[26] | proc_34_data_PIPO_blk[26] | proc_34_start_FIFO_blk[26] | proc_34_TLF_FIFO_blk[26] | proc_34_input_sync_blk[26] | proc_34_output_sync_blk[26]);
    assign proc_34_data_FIFO_blk[27] = 1'b0;
    assign proc_34_data_PIPO_blk[27] = 1'b0;
    assign proc_34_start_FIFO_blk[27] = 1'b0;
    assign proc_34_TLF_FIFO_blk[27] = 1'b0;
    assign proc_34_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_34_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_34[27] = dl_detect_out ? proc_dep_vld_vec_34_reg[27] : (proc_34_data_FIFO_blk[27] | proc_34_data_PIPO_blk[27] | proc_34_start_FIFO_blk[27] | proc_34_TLF_FIFO_blk[27] | proc_34_input_sync_blk[27] | proc_34_output_sync_blk[27]);
    assign proc_34_data_FIFO_blk[28] = 1'b0;
    assign proc_34_data_PIPO_blk[28] = 1'b0;
    assign proc_34_start_FIFO_blk[28] = 1'b0;
    assign proc_34_TLF_FIFO_blk[28] = 1'b0;
    assign proc_34_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_34_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_34[28] = dl_detect_out ? proc_dep_vld_vec_34_reg[28] : (proc_34_data_FIFO_blk[28] | proc_34_data_PIPO_blk[28] | proc_34_start_FIFO_blk[28] | proc_34_TLF_FIFO_blk[28] | proc_34_input_sync_blk[28] | proc_34_output_sync_blk[28]);
    assign proc_34_data_FIFO_blk[29] = 1'b0;
    assign proc_34_data_PIPO_blk[29] = 1'b0;
    assign proc_34_start_FIFO_blk[29] = 1'b0;
    assign proc_34_TLF_FIFO_blk[29] = 1'b0;
    assign proc_34_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_34_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_34[29] = dl_detect_out ? proc_dep_vld_vec_34_reg[29] : (proc_34_data_FIFO_blk[29] | proc_34_data_PIPO_blk[29] | proc_34_start_FIFO_blk[29] | proc_34_TLF_FIFO_blk[29] | proc_34_input_sync_blk[29] | proc_34_output_sync_blk[29]);
    assign proc_34_data_FIFO_blk[30] = 1'b0;
    assign proc_34_data_PIPO_blk[30] = 1'b0;
    assign proc_34_start_FIFO_blk[30] = 1'b0;
    assign proc_34_TLF_FIFO_blk[30] = 1'b0;
    assign proc_34_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_34_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_34[30] = dl_detect_out ? proc_dep_vld_vec_34_reg[30] : (proc_34_data_FIFO_blk[30] | proc_34_data_PIPO_blk[30] | proc_34_start_FIFO_blk[30] | proc_34_TLF_FIFO_blk[30] | proc_34_input_sync_blk[30] | proc_34_output_sync_blk[30]);
    assign proc_34_data_FIFO_blk[31] = 1'b0;
    assign proc_34_data_PIPO_blk[31] = 1'b0;
    assign proc_34_start_FIFO_blk[31] = 1'b0;
    assign proc_34_TLF_FIFO_blk[31] = 1'b0;
    assign proc_34_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_34_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_34[31] = dl_detect_out ? proc_dep_vld_vec_34_reg[31] : (proc_34_data_FIFO_blk[31] | proc_34_data_PIPO_blk[31] | proc_34_start_FIFO_blk[31] | proc_34_TLF_FIFO_blk[31] | proc_34_input_sync_blk[31] | proc_34_output_sync_blk[31]);
    assign proc_34_data_FIFO_blk[32] = 1'b0;
    assign proc_34_data_PIPO_blk[32] = 1'b0;
    assign proc_34_start_FIFO_blk[32] = 1'b0;
    assign proc_34_TLF_FIFO_blk[32] = 1'b0;
    assign proc_34_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_29_U0_ap_ready & ProcessingElement_29_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_34_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_34[32] = dl_detect_out ? proc_dep_vld_vec_34_reg[32] : (proc_34_data_FIFO_blk[32] | proc_34_data_PIPO_blk[32] | proc_34_start_FIFO_blk[32] | proc_34_TLF_FIFO_blk[32] | proc_34_input_sync_blk[32] | proc_34_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_34_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_34_reg <= proc_dep_vld_vec_34;
        end
    end
    assign in_chan_dep_vld_vec_34[0] = dep_chan_vld_0_34;
    assign in_chan_dep_data_vec_34[39 : 0] = dep_chan_data_0_34;
    assign token_in_vec_34[0] = token_0_34;
    assign in_chan_dep_vld_vec_34[1] = dep_chan_vld_1_34;
    assign in_chan_dep_data_vec_34[79 : 40] = dep_chan_data_1_34;
    assign token_in_vec_34[1] = token_1_34;
    assign in_chan_dep_vld_vec_34[2] = dep_chan_vld_3_34;
    assign in_chan_dep_data_vec_34[119 : 80] = dep_chan_data_3_34;
    assign token_in_vec_34[2] = token_3_34;
    assign in_chan_dep_vld_vec_34[3] = dep_chan_vld_6_34;
    assign in_chan_dep_data_vec_34[159 : 120] = dep_chan_data_6_34;
    assign token_in_vec_34[3] = token_6_34;
    assign in_chan_dep_vld_vec_34[4] = dep_chan_vld_7_34;
    assign in_chan_dep_data_vec_34[199 : 160] = dep_chan_data_7_34;
    assign token_in_vec_34[4] = token_7_34;
    assign in_chan_dep_vld_vec_34[5] = dep_chan_vld_8_34;
    assign in_chan_dep_data_vec_34[239 : 200] = dep_chan_data_8_34;
    assign token_in_vec_34[5] = token_8_34;
    assign in_chan_dep_vld_vec_34[6] = dep_chan_vld_9_34;
    assign in_chan_dep_data_vec_34[279 : 240] = dep_chan_data_9_34;
    assign token_in_vec_34[6] = token_9_34;
    assign in_chan_dep_vld_vec_34[7] = dep_chan_vld_10_34;
    assign in_chan_dep_data_vec_34[319 : 280] = dep_chan_data_10_34;
    assign token_in_vec_34[7] = token_10_34;
    assign in_chan_dep_vld_vec_34[8] = dep_chan_vld_11_34;
    assign in_chan_dep_data_vec_34[359 : 320] = dep_chan_data_11_34;
    assign token_in_vec_34[8] = token_11_34;
    assign in_chan_dep_vld_vec_34[9] = dep_chan_vld_12_34;
    assign in_chan_dep_data_vec_34[399 : 360] = dep_chan_data_12_34;
    assign token_in_vec_34[9] = token_12_34;
    assign in_chan_dep_vld_vec_34[10] = dep_chan_vld_13_34;
    assign in_chan_dep_data_vec_34[439 : 400] = dep_chan_data_13_34;
    assign token_in_vec_34[10] = token_13_34;
    assign in_chan_dep_vld_vec_34[11] = dep_chan_vld_14_34;
    assign in_chan_dep_data_vec_34[479 : 440] = dep_chan_data_14_34;
    assign token_in_vec_34[11] = token_14_34;
    assign in_chan_dep_vld_vec_34[12] = dep_chan_vld_15_34;
    assign in_chan_dep_data_vec_34[519 : 480] = dep_chan_data_15_34;
    assign token_in_vec_34[12] = token_15_34;
    assign in_chan_dep_vld_vec_34[13] = dep_chan_vld_16_34;
    assign in_chan_dep_data_vec_34[559 : 520] = dep_chan_data_16_34;
    assign token_in_vec_34[13] = token_16_34;
    assign in_chan_dep_vld_vec_34[14] = dep_chan_vld_17_34;
    assign in_chan_dep_data_vec_34[599 : 560] = dep_chan_data_17_34;
    assign token_in_vec_34[14] = token_17_34;
    assign in_chan_dep_vld_vec_34[15] = dep_chan_vld_18_34;
    assign in_chan_dep_data_vec_34[639 : 600] = dep_chan_data_18_34;
    assign token_in_vec_34[15] = token_18_34;
    assign in_chan_dep_vld_vec_34[16] = dep_chan_vld_19_34;
    assign in_chan_dep_data_vec_34[679 : 640] = dep_chan_data_19_34;
    assign token_in_vec_34[16] = token_19_34;
    assign in_chan_dep_vld_vec_34[17] = dep_chan_vld_20_34;
    assign in_chan_dep_data_vec_34[719 : 680] = dep_chan_data_20_34;
    assign token_in_vec_34[17] = token_20_34;
    assign in_chan_dep_vld_vec_34[18] = dep_chan_vld_21_34;
    assign in_chan_dep_data_vec_34[759 : 720] = dep_chan_data_21_34;
    assign token_in_vec_34[18] = token_21_34;
    assign in_chan_dep_vld_vec_34[19] = dep_chan_vld_22_34;
    assign in_chan_dep_data_vec_34[799 : 760] = dep_chan_data_22_34;
    assign token_in_vec_34[19] = token_22_34;
    assign in_chan_dep_vld_vec_34[20] = dep_chan_vld_23_34;
    assign in_chan_dep_data_vec_34[839 : 800] = dep_chan_data_23_34;
    assign token_in_vec_34[20] = token_23_34;
    assign in_chan_dep_vld_vec_34[21] = dep_chan_vld_24_34;
    assign in_chan_dep_data_vec_34[879 : 840] = dep_chan_data_24_34;
    assign token_in_vec_34[21] = token_24_34;
    assign in_chan_dep_vld_vec_34[22] = dep_chan_vld_25_34;
    assign in_chan_dep_data_vec_34[919 : 880] = dep_chan_data_25_34;
    assign token_in_vec_34[22] = token_25_34;
    assign in_chan_dep_vld_vec_34[23] = dep_chan_vld_26_34;
    assign in_chan_dep_data_vec_34[959 : 920] = dep_chan_data_26_34;
    assign token_in_vec_34[23] = token_26_34;
    assign in_chan_dep_vld_vec_34[24] = dep_chan_vld_27_34;
    assign in_chan_dep_data_vec_34[999 : 960] = dep_chan_data_27_34;
    assign token_in_vec_34[24] = token_27_34;
    assign in_chan_dep_vld_vec_34[25] = dep_chan_vld_28_34;
    assign in_chan_dep_data_vec_34[1039 : 1000] = dep_chan_data_28_34;
    assign token_in_vec_34[25] = token_28_34;
    assign in_chan_dep_vld_vec_34[26] = dep_chan_vld_29_34;
    assign in_chan_dep_data_vec_34[1079 : 1040] = dep_chan_data_29_34;
    assign token_in_vec_34[26] = token_29_34;
    assign in_chan_dep_vld_vec_34[27] = dep_chan_vld_30_34;
    assign in_chan_dep_data_vec_34[1119 : 1080] = dep_chan_data_30_34;
    assign token_in_vec_34[27] = token_30_34;
    assign in_chan_dep_vld_vec_34[28] = dep_chan_vld_31_34;
    assign in_chan_dep_data_vec_34[1159 : 1120] = dep_chan_data_31_34;
    assign token_in_vec_34[28] = token_31_34;
    assign in_chan_dep_vld_vec_34[29] = dep_chan_vld_32_34;
    assign in_chan_dep_data_vec_34[1199 : 1160] = dep_chan_data_32_34;
    assign token_in_vec_34[29] = token_32_34;
    assign in_chan_dep_vld_vec_34[30] = dep_chan_vld_33_34;
    assign in_chan_dep_data_vec_34[1239 : 1200] = dep_chan_data_33_34;
    assign token_in_vec_34[30] = token_33_34;
    assign in_chan_dep_vld_vec_34[31] = dep_chan_vld_35_34;
    assign in_chan_dep_data_vec_34[1279 : 1240] = dep_chan_data_35_34;
    assign token_in_vec_34[31] = token_35_34;
    assign in_chan_dep_vld_vec_34[32] = dep_chan_vld_36_34;
    assign in_chan_dep_data_vec_34[1319 : 1280] = dep_chan_data_36_34;
    assign token_in_vec_34[32] = token_36_34;
    assign dep_chan_vld_34_33 = out_chan_dep_vld_vec_34[0];
    assign dep_chan_data_34_33 = out_chan_dep_data_34;
    assign token_34_33 = token_out_vec_34[0];
    assign dep_chan_vld_34_35 = out_chan_dep_vld_vec_34[1];
    assign dep_chan_data_34_35 = out_chan_dep_data_34;
    assign token_34_35 = token_out_vec_34[1];
    assign dep_chan_vld_34_0 = out_chan_dep_vld_vec_34[2];
    assign dep_chan_data_34_0 = out_chan_dep_data_34;
    assign token_34_0 = token_out_vec_34[2];
    assign dep_chan_vld_34_1 = out_chan_dep_vld_vec_34[3];
    assign dep_chan_data_34_1 = out_chan_dep_data_34;
    assign token_34_1 = token_out_vec_34[3];
    assign dep_chan_vld_34_3 = out_chan_dep_vld_vec_34[4];
    assign dep_chan_data_34_3 = out_chan_dep_data_34;
    assign token_34_3 = token_out_vec_34[4];
    assign dep_chan_vld_34_6 = out_chan_dep_vld_vec_34[5];
    assign dep_chan_data_34_6 = out_chan_dep_data_34;
    assign token_34_6 = token_out_vec_34[5];
    assign dep_chan_vld_34_7 = out_chan_dep_vld_vec_34[6];
    assign dep_chan_data_34_7 = out_chan_dep_data_34;
    assign token_34_7 = token_out_vec_34[6];
    assign dep_chan_vld_34_8 = out_chan_dep_vld_vec_34[7];
    assign dep_chan_data_34_8 = out_chan_dep_data_34;
    assign token_34_8 = token_out_vec_34[7];
    assign dep_chan_vld_34_9 = out_chan_dep_vld_vec_34[8];
    assign dep_chan_data_34_9 = out_chan_dep_data_34;
    assign token_34_9 = token_out_vec_34[8];
    assign dep_chan_vld_34_10 = out_chan_dep_vld_vec_34[9];
    assign dep_chan_data_34_10 = out_chan_dep_data_34;
    assign token_34_10 = token_out_vec_34[9];
    assign dep_chan_vld_34_11 = out_chan_dep_vld_vec_34[10];
    assign dep_chan_data_34_11 = out_chan_dep_data_34;
    assign token_34_11 = token_out_vec_34[10];
    assign dep_chan_vld_34_12 = out_chan_dep_vld_vec_34[11];
    assign dep_chan_data_34_12 = out_chan_dep_data_34;
    assign token_34_12 = token_out_vec_34[11];
    assign dep_chan_vld_34_13 = out_chan_dep_vld_vec_34[12];
    assign dep_chan_data_34_13 = out_chan_dep_data_34;
    assign token_34_13 = token_out_vec_34[12];
    assign dep_chan_vld_34_14 = out_chan_dep_vld_vec_34[13];
    assign dep_chan_data_34_14 = out_chan_dep_data_34;
    assign token_34_14 = token_out_vec_34[13];
    assign dep_chan_vld_34_15 = out_chan_dep_vld_vec_34[14];
    assign dep_chan_data_34_15 = out_chan_dep_data_34;
    assign token_34_15 = token_out_vec_34[14];
    assign dep_chan_vld_34_16 = out_chan_dep_vld_vec_34[15];
    assign dep_chan_data_34_16 = out_chan_dep_data_34;
    assign token_34_16 = token_out_vec_34[15];
    assign dep_chan_vld_34_17 = out_chan_dep_vld_vec_34[16];
    assign dep_chan_data_34_17 = out_chan_dep_data_34;
    assign token_34_17 = token_out_vec_34[16];
    assign dep_chan_vld_34_18 = out_chan_dep_vld_vec_34[17];
    assign dep_chan_data_34_18 = out_chan_dep_data_34;
    assign token_34_18 = token_out_vec_34[17];
    assign dep_chan_vld_34_19 = out_chan_dep_vld_vec_34[18];
    assign dep_chan_data_34_19 = out_chan_dep_data_34;
    assign token_34_19 = token_out_vec_34[18];
    assign dep_chan_vld_34_20 = out_chan_dep_vld_vec_34[19];
    assign dep_chan_data_34_20 = out_chan_dep_data_34;
    assign token_34_20 = token_out_vec_34[19];
    assign dep_chan_vld_34_21 = out_chan_dep_vld_vec_34[20];
    assign dep_chan_data_34_21 = out_chan_dep_data_34;
    assign token_34_21 = token_out_vec_34[20];
    assign dep_chan_vld_34_22 = out_chan_dep_vld_vec_34[21];
    assign dep_chan_data_34_22 = out_chan_dep_data_34;
    assign token_34_22 = token_out_vec_34[21];
    assign dep_chan_vld_34_23 = out_chan_dep_vld_vec_34[22];
    assign dep_chan_data_34_23 = out_chan_dep_data_34;
    assign token_34_23 = token_out_vec_34[22];
    assign dep_chan_vld_34_24 = out_chan_dep_vld_vec_34[23];
    assign dep_chan_data_34_24 = out_chan_dep_data_34;
    assign token_34_24 = token_out_vec_34[23];
    assign dep_chan_vld_34_25 = out_chan_dep_vld_vec_34[24];
    assign dep_chan_data_34_25 = out_chan_dep_data_34;
    assign token_34_25 = token_out_vec_34[24];
    assign dep_chan_vld_34_26 = out_chan_dep_vld_vec_34[25];
    assign dep_chan_data_34_26 = out_chan_dep_data_34;
    assign token_34_26 = token_out_vec_34[25];
    assign dep_chan_vld_34_27 = out_chan_dep_vld_vec_34[26];
    assign dep_chan_data_34_27 = out_chan_dep_data_34;
    assign token_34_27 = token_out_vec_34[26];
    assign dep_chan_vld_34_28 = out_chan_dep_vld_vec_34[27];
    assign dep_chan_data_34_28 = out_chan_dep_data_34;
    assign token_34_28 = token_out_vec_34[27];
    assign dep_chan_vld_34_29 = out_chan_dep_vld_vec_34[28];
    assign dep_chan_data_34_29 = out_chan_dep_data_34;
    assign token_34_29 = token_out_vec_34[28];
    assign dep_chan_vld_34_30 = out_chan_dep_vld_vec_34[29];
    assign dep_chan_data_34_30 = out_chan_dep_data_34;
    assign token_34_30 = token_out_vec_34[29];
    assign dep_chan_vld_34_31 = out_chan_dep_vld_vec_34[30];
    assign dep_chan_data_34_31 = out_chan_dep_data_34;
    assign token_34_31 = token_out_vec_34[30];
    assign dep_chan_vld_34_32 = out_chan_dep_vld_vec_34[31];
    assign dep_chan_data_34_32 = out_chan_dep_data_34;
    assign token_34_32 = token_out_vec_34[31];
    assign dep_chan_vld_34_36 = out_chan_dep_vld_vec_34[32];
    assign dep_chan_data_34_36 = out_chan_dep_data_34;
    assign token_34_36 = token_out_vec_34[32];

    // Process: ProcessingElement_30_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 35, 33, 33) MatrixMultiplicationKernel_hls_deadlock_detect_unit_35 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_35),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_35),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_35),
        .token_in_vec(token_in_vec_35),
        .dl_detect_in(dl_detect_out),
        .origin(origin[35]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_35),
        .out_chan_dep_data(out_chan_dep_data_35),
        .token_out_vec(token_out_vec_35),
        .dl_detect_out(dl_in_vec[35]));

    assign proc_35_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_29_blk_n) | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_29_blk_n) | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_WriteC_Flattened_fu_179.cPipes_29_blk_n);
    assign proc_35_data_PIPO_blk[0] = 1'b0;
    assign proc_35_start_FIFO_blk[0] = 1'b0;
    assign proc_35_TLF_FIFO_blk[0] = 1'b0;
    assign proc_35_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_35_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_35[0] = dl_detect_out ? proc_dep_vld_vec_35_reg[0] : (proc_35_data_FIFO_blk[0] | proc_35_data_PIPO_blk[0] | proc_35_start_FIFO_blk[0] | proc_35_TLF_FIFO_blk[0] | proc_35_input_sync_blk[0] | proc_35_output_sync_blk[0]);
    assign proc_35_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_Pipeline_N_Pipeline_M_fu_157.aPipes_30_blk_n) | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_Pipeline_N_Pipeline_M_fu_157.bPipes_30_blk_n) | (~ProcessingElement_30_U0.grp_ProcessingElement_30_Pipeline_WriteC_Flattened_fu_179.cPipes_30_blk_n);
    assign proc_35_data_PIPO_blk[1] = 1'b0;
    assign proc_35_start_FIFO_blk[1] = 1'b0;
    assign proc_35_TLF_FIFO_blk[1] = 1'b0;
    assign proc_35_input_sync_blk[1] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_31_U0_ap_ready);
    assign proc_35_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_35[1] = dl_detect_out ? proc_dep_vld_vec_35_reg[1] : (proc_35_data_FIFO_blk[1] | proc_35_data_PIPO_blk[1] | proc_35_start_FIFO_blk[1] | proc_35_TLF_FIFO_blk[1] | proc_35_input_sync_blk[1] | proc_35_output_sync_blk[1]);
    assign proc_35_data_FIFO_blk[2] = 1'b0;
    assign proc_35_data_PIPO_blk[2] = 1'b0;
    assign proc_35_start_FIFO_blk[2] = 1'b0;
    assign proc_35_TLF_FIFO_blk[2] = 1'b0;
    assign proc_35_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_35_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_35[2] = dl_detect_out ? proc_dep_vld_vec_35_reg[2] : (proc_35_data_FIFO_blk[2] | proc_35_data_PIPO_blk[2] | proc_35_start_FIFO_blk[2] | proc_35_TLF_FIFO_blk[2] | proc_35_input_sync_blk[2] | proc_35_output_sync_blk[2]);
    assign proc_35_data_FIFO_blk[3] = 1'b0;
    assign proc_35_data_PIPO_blk[3] = 1'b0;
    assign proc_35_start_FIFO_blk[3] = 1'b0;
    assign proc_35_TLF_FIFO_blk[3] = 1'b0;
    assign proc_35_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_35_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_35[3] = dl_detect_out ? proc_dep_vld_vec_35_reg[3] : (proc_35_data_FIFO_blk[3] | proc_35_data_PIPO_blk[3] | proc_35_start_FIFO_blk[3] | proc_35_TLF_FIFO_blk[3] | proc_35_input_sync_blk[3] | proc_35_output_sync_blk[3]);
    assign proc_35_data_FIFO_blk[4] = 1'b0;
    assign proc_35_data_PIPO_blk[4] = 1'b0;
    assign proc_35_start_FIFO_blk[4] = 1'b0;
    assign proc_35_TLF_FIFO_blk[4] = 1'b0;
    assign proc_35_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_35_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_35[4] = dl_detect_out ? proc_dep_vld_vec_35_reg[4] : (proc_35_data_FIFO_blk[4] | proc_35_data_PIPO_blk[4] | proc_35_start_FIFO_blk[4] | proc_35_TLF_FIFO_blk[4] | proc_35_input_sync_blk[4] | proc_35_output_sync_blk[4]);
    assign proc_35_data_FIFO_blk[5] = 1'b0;
    assign proc_35_data_PIPO_blk[5] = 1'b0;
    assign proc_35_start_FIFO_blk[5] = 1'b0;
    assign proc_35_TLF_FIFO_blk[5] = 1'b0;
    assign proc_35_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_35_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_35[5] = dl_detect_out ? proc_dep_vld_vec_35_reg[5] : (proc_35_data_FIFO_blk[5] | proc_35_data_PIPO_blk[5] | proc_35_start_FIFO_blk[5] | proc_35_TLF_FIFO_blk[5] | proc_35_input_sync_blk[5] | proc_35_output_sync_blk[5]);
    assign proc_35_data_FIFO_blk[6] = 1'b0;
    assign proc_35_data_PIPO_blk[6] = 1'b0;
    assign proc_35_start_FIFO_blk[6] = 1'b0;
    assign proc_35_TLF_FIFO_blk[6] = 1'b0;
    assign proc_35_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_35_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_35[6] = dl_detect_out ? proc_dep_vld_vec_35_reg[6] : (proc_35_data_FIFO_blk[6] | proc_35_data_PIPO_blk[6] | proc_35_start_FIFO_blk[6] | proc_35_TLF_FIFO_blk[6] | proc_35_input_sync_blk[6] | proc_35_output_sync_blk[6]);
    assign proc_35_data_FIFO_blk[7] = 1'b0;
    assign proc_35_data_PIPO_blk[7] = 1'b0;
    assign proc_35_start_FIFO_blk[7] = 1'b0;
    assign proc_35_TLF_FIFO_blk[7] = 1'b0;
    assign proc_35_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_35_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_35[7] = dl_detect_out ? proc_dep_vld_vec_35_reg[7] : (proc_35_data_FIFO_blk[7] | proc_35_data_PIPO_blk[7] | proc_35_start_FIFO_blk[7] | proc_35_TLF_FIFO_blk[7] | proc_35_input_sync_blk[7] | proc_35_output_sync_blk[7]);
    assign proc_35_data_FIFO_blk[8] = 1'b0;
    assign proc_35_data_PIPO_blk[8] = 1'b0;
    assign proc_35_start_FIFO_blk[8] = 1'b0;
    assign proc_35_TLF_FIFO_blk[8] = 1'b0;
    assign proc_35_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_35_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_35[8] = dl_detect_out ? proc_dep_vld_vec_35_reg[8] : (proc_35_data_FIFO_blk[8] | proc_35_data_PIPO_blk[8] | proc_35_start_FIFO_blk[8] | proc_35_TLF_FIFO_blk[8] | proc_35_input_sync_blk[8] | proc_35_output_sync_blk[8]);
    assign proc_35_data_FIFO_blk[9] = 1'b0;
    assign proc_35_data_PIPO_blk[9] = 1'b0;
    assign proc_35_start_FIFO_blk[9] = 1'b0;
    assign proc_35_TLF_FIFO_blk[9] = 1'b0;
    assign proc_35_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_35_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_35[9] = dl_detect_out ? proc_dep_vld_vec_35_reg[9] : (proc_35_data_FIFO_blk[9] | proc_35_data_PIPO_blk[9] | proc_35_start_FIFO_blk[9] | proc_35_TLF_FIFO_blk[9] | proc_35_input_sync_blk[9] | proc_35_output_sync_blk[9]);
    assign proc_35_data_FIFO_blk[10] = 1'b0;
    assign proc_35_data_PIPO_blk[10] = 1'b0;
    assign proc_35_start_FIFO_blk[10] = 1'b0;
    assign proc_35_TLF_FIFO_blk[10] = 1'b0;
    assign proc_35_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_35_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_35[10] = dl_detect_out ? proc_dep_vld_vec_35_reg[10] : (proc_35_data_FIFO_blk[10] | proc_35_data_PIPO_blk[10] | proc_35_start_FIFO_blk[10] | proc_35_TLF_FIFO_blk[10] | proc_35_input_sync_blk[10] | proc_35_output_sync_blk[10]);
    assign proc_35_data_FIFO_blk[11] = 1'b0;
    assign proc_35_data_PIPO_blk[11] = 1'b0;
    assign proc_35_start_FIFO_blk[11] = 1'b0;
    assign proc_35_TLF_FIFO_blk[11] = 1'b0;
    assign proc_35_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_35_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_35[11] = dl_detect_out ? proc_dep_vld_vec_35_reg[11] : (proc_35_data_FIFO_blk[11] | proc_35_data_PIPO_blk[11] | proc_35_start_FIFO_blk[11] | proc_35_TLF_FIFO_blk[11] | proc_35_input_sync_blk[11] | proc_35_output_sync_blk[11]);
    assign proc_35_data_FIFO_blk[12] = 1'b0;
    assign proc_35_data_PIPO_blk[12] = 1'b0;
    assign proc_35_start_FIFO_blk[12] = 1'b0;
    assign proc_35_TLF_FIFO_blk[12] = 1'b0;
    assign proc_35_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_35_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_35[12] = dl_detect_out ? proc_dep_vld_vec_35_reg[12] : (proc_35_data_FIFO_blk[12] | proc_35_data_PIPO_blk[12] | proc_35_start_FIFO_blk[12] | proc_35_TLF_FIFO_blk[12] | proc_35_input_sync_blk[12] | proc_35_output_sync_blk[12]);
    assign proc_35_data_FIFO_blk[13] = 1'b0;
    assign proc_35_data_PIPO_blk[13] = 1'b0;
    assign proc_35_start_FIFO_blk[13] = 1'b0;
    assign proc_35_TLF_FIFO_blk[13] = 1'b0;
    assign proc_35_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_35_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_35[13] = dl_detect_out ? proc_dep_vld_vec_35_reg[13] : (proc_35_data_FIFO_blk[13] | proc_35_data_PIPO_blk[13] | proc_35_start_FIFO_blk[13] | proc_35_TLF_FIFO_blk[13] | proc_35_input_sync_blk[13] | proc_35_output_sync_blk[13]);
    assign proc_35_data_FIFO_blk[14] = 1'b0;
    assign proc_35_data_PIPO_blk[14] = 1'b0;
    assign proc_35_start_FIFO_blk[14] = 1'b0;
    assign proc_35_TLF_FIFO_blk[14] = 1'b0;
    assign proc_35_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_35_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_35[14] = dl_detect_out ? proc_dep_vld_vec_35_reg[14] : (proc_35_data_FIFO_blk[14] | proc_35_data_PIPO_blk[14] | proc_35_start_FIFO_blk[14] | proc_35_TLF_FIFO_blk[14] | proc_35_input_sync_blk[14] | proc_35_output_sync_blk[14]);
    assign proc_35_data_FIFO_blk[15] = 1'b0;
    assign proc_35_data_PIPO_blk[15] = 1'b0;
    assign proc_35_start_FIFO_blk[15] = 1'b0;
    assign proc_35_TLF_FIFO_blk[15] = 1'b0;
    assign proc_35_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_35_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_35[15] = dl_detect_out ? proc_dep_vld_vec_35_reg[15] : (proc_35_data_FIFO_blk[15] | proc_35_data_PIPO_blk[15] | proc_35_start_FIFO_blk[15] | proc_35_TLF_FIFO_blk[15] | proc_35_input_sync_blk[15] | proc_35_output_sync_blk[15]);
    assign proc_35_data_FIFO_blk[16] = 1'b0;
    assign proc_35_data_PIPO_blk[16] = 1'b0;
    assign proc_35_start_FIFO_blk[16] = 1'b0;
    assign proc_35_TLF_FIFO_blk[16] = 1'b0;
    assign proc_35_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_35_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_35[16] = dl_detect_out ? proc_dep_vld_vec_35_reg[16] : (proc_35_data_FIFO_blk[16] | proc_35_data_PIPO_blk[16] | proc_35_start_FIFO_blk[16] | proc_35_TLF_FIFO_blk[16] | proc_35_input_sync_blk[16] | proc_35_output_sync_blk[16]);
    assign proc_35_data_FIFO_blk[17] = 1'b0;
    assign proc_35_data_PIPO_blk[17] = 1'b0;
    assign proc_35_start_FIFO_blk[17] = 1'b0;
    assign proc_35_TLF_FIFO_blk[17] = 1'b0;
    assign proc_35_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_35_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_35[17] = dl_detect_out ? proc_dep_vld_vec_35_reg[17] : (proc_35_data_FIFO_blk[17] | proc_35_data_PIPO_blk[17] | proc_35_start_FIFO_blk[17] | proc_35_TLF_FIFO_blk[17] | proc_35_input_sync_blk[17] | proc_35_output_sync_blk[17]);
    assign proc_35_data_FIFO_blk[18] = 1'b0;
    assign proc_35_data_PIPO_blk[18] = 1'b0;
    assign proc_35_start_FIFO_blk[18] = 1'b0;
    assign proc_35_TLF_FIFO_blk[18] = 1'b0;
    assign proc_35_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_35_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_35[18] = dl_detect_out ? proc_dep_vld_vec_35_reg[18] : (proc_35_data_FIFO_blk[18] | proc_35_data_PIPO_blk[18] | proc_35_start_FIFO_blk[18] | proc_35_TLF_FIFO_blk[18] | proc_35_input_sync_blk[18] | proc_35_output_sync_blk[18]);
    assign proc_35_data_FIFO_blk[19] = 1'b0;
    assign proc_35_data_PIPO_blk[19] = 1'b0;
    assign proc_35_start_FIFO_blk[19] = 1'b0;
    assign proc_35_TLF_FIFO_blk[19] = 1'b0;
    assign proc_35_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_35_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_35[19] = dl_detect_out ? proc_dep_vld_vec_35_reg[19] : (proc_35_data_FIFO_blk[19] | proc_35_data_PIPO_blk[19] | proc_35_start_FIFO_blk[19] | proc_35_TLF_FIFO_blk[19] | proc_35_input_sync_blk[19] | proc_35_output_sync_blk[19]);
    assign proc_35_data_FIFO_blk[20] = 1'b0;
    assign proc_35_data_PIPO_blk[20] = 1'b0;
    assign proc_35_start_FIFO_blk[20] = 1'b0;
    assign proc_35_TLF_FIFO_blk[20] = 1'b0;
    assign proc_35_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_35_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_35[20] = dl_detect_out ? proc_dep_vld_vec_35_reg[20] : (proc_35_data_FIFO_blk[20] | proc_35_data_PIPO_blk[20] | proc_35_start_FIFO_blk[20] | proc_35_TLF_FIFO_blk[20] | proc_35_input_sync_blk[20] | proc_35_output_sync_blk[20]);
    assign proc_35_data_FIFO_blk[21] = 1'b0;
    assign proc_35_data_PIPO_blk[21] = 1'b0;
    assign proc_35_start_FIFO_blk[21] = 1'b0;
    assign proc_35_TLF_FIFO_blk[21] = 1'b0;
    assign proc_35_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_35_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_35[21] = dl_detect_out ? proc_dep_vld_vec_35_reg[21] : (proc_35_data_FIFO_blk[21] | proc_35_data_PIPO_blk[21] | proc_35_start_FIFO_blk[21] | proc_35_TLF_FIFO_blk[21] | proc_35_input_sync_blk[21] | proc_35_output_sync_blk[21]);
    assign proc_35_data_FIFO_blk[22] = 1'b0;
    assign proc_35_data_PIPO_blk[22] = 1'b0;
    assign proc_35_start_FIFO_blk[22] = 1'b0;
    assign proc_35_TLF_FIFO_blk[22] = 1'b0;
    assign proc_35_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_35_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_35[22] = dl_detect_out ? proc_dep_vld_vec_35_reg[22] : (proc_35_data_FIFO_blk[22] | proc_35_data_PIPO_blk[22] | proc_35_start_FIFO_blk[22] | proc_35_TLF_FIFO_blk[22] | proc_35_input_sync_blk[22] | proc_35_output_sync_blk[22]);
    assign proc_35_data_FIFO_blk[23] = 1'b0;
    assign proc_35_data_PIPO_blk[23] = 1'b0;
    assign proc_35_start_FIFO_blk[23] = 1'b0;
    assign proc_35_TLF_FIFO_blk[23] = 1'b0;
    assign proc_35_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_35_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_35[23] = dl_detect_out ? proc_dep_vld_vec_35_reg[23] : (proc_35_data_FIFO_blk[23] | proc_35_data_PIPO_blk[23] | proc_35_start_FIFO_blk[23] | proc_35_TLF_FIFO_blk[23] | proc_35_input_sync_blk[23] | proc_35_output_sync_blk[23]);
    assign proc_35_data_FIFO_blk[24] = 1'b0;
    assign proc_35_data_PIPO_blk[24] = 1'b0;
    assign proc_35_start_FIFO_blk[24] = 1'b0;
    assign proc_35_TLF_FIFO_blk[24] = 1'b0;
    assign proc_35_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_35_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_35[24] = dl_detect_out ? proc_dep_vld_vec_35_reg[24] : (proc_35_data_FIFO_blk[24] | proc_35_data_PIPO_blk[24] | proc_35_start_FIFO_blk[24] | proc_35_TLF_FIFO_blk[24] | proc_35_input_sync_blk[24] | proc_35_output_sync_blk[24]);
    assign proc_35_data_FIFO_blk[25] = 1'b0;
    assign proc_35_data_PIPO_blk[25] = 1'b0;
    assign proc_35_start_FIFO_blk[25] = 1'b0;
    assign proc_35_TLF_FIFO_blk[25] = 1'b0;
    assign proc_35_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_35_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_35[25] = dl_detect_out ? proc_dep_vld_vec_35_reg[25] : (proc_35_data_FIFO_blk[25] | proc_35_data_PIPO_blk[25] | proc_35_start_FIFO_blk[25] | proc_35_TLF_FIFO_blk[25] | proc_35_input_sync_blk[25] | proc_35_output_sync_blk[25]);
    assign proc_35_data_FIFO_blk[26] = 1'b0;
    assign proc_35_data_PIPO_blk[26] = 1'b0;
    assign proc_35_start_FIFO_blk[26] = 1'b0;
    assign proc_35_TLF_FIFO_blk[26] = 1'b0;
    assign proc_35_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_35_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_35[26] = dl_detect_out ? proc_dep_vld_vec_35_reg[26] : (proc_35_data_FIFO_blk[26] | proc_35_data_PIPO_blk[26] | proc_35_start_FIFO_blk[26] | proc_35_TLF_FIFO_blk[26] | proc_35_input_sync_blk[26] | proc_35_output_sync_blk[26]);
    assign proc_35_data_FIFO_blk[27] = 1'b0;
    assign proc_35_data_PIPO_blk[27] = 1'b0;
    assign proc_35_start_FIFO_blk[27] = 1'b0;
    assign proc_35_TLF_FIFO_blk[27] = 1'b0;
    assign proc_35_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_35_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_35[27] = dl_detect_out ? proc_dep_vld_vec_35_reg[27] : (proc_35_data_FIFO_blk[27] | proc_35_data_PIPO_blk[27] | proc_35_start_FIFO_blk[27] | proc_35_TLF_FIFO_blk[27] | proc_35_input_sync_blk[27] | proc_35_output_sync_blk[27]);
    assign proc_35_data_FIFO_blk[28] = 1'b0;
    assign proc_35_data_PIPO_blk[28] = 1'b0;
    assign proc_35_start_FIFO_blk[28] = 1'b0;
    assign proc_35_TLF_FIFO_blk[28] = 1'b0;
    assign proc_35_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_35_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_35[28] = dl_detect_out ? proc_dep_vld_vec_35_reg[28] : (proc_35_data_FIFO_blk[28] | proc_35_data_PIPO_blk[28] | proc_35_start_FIFO_blk[28] | proc_35_TLF_FIFO_blk[28] | proc_35_input_sync_blk[28] | proc_35_output_sync_blk[28]);
    assign proc_35_data_FIFO_blk[29] = 1'b0;
    assign proc_35_data_PIPO_blk[29] = 1'b0;
    assign proc_35_start_FIFO_blk[29] = 1'b0;
    assign proc_35_TLF_FIFO_blk[29] = 1'b0;
    assign proc_35_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_35_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_35[29] = dl_detect_out ? proc_dep_vld_vec_35_reg[29] : (proc_35_data_FIFO_blk[29] | proc_35_data_PIPO_blk[29] | proc_35_start_FIFO_blk[29] | proc_35_TLF_FIFO_blk[29] | proc_35_input_sync_blk[29] | proc_35_output_sync_blk[29]);
    assign proc_35_data_FIFO_blk[30] = 1'b0;
    assign proc_35_data_PIPO_blk[30] = 1'b0;
    assign proc_35_start_FIFO_blk[30] = 1'b0;
    assign proc_35_TLF_FIFO_blk[30] = 1'b0;
    assign proc_35_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_35_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_35[30] = dl_detect_out ? proc_dep_vld_vec_35_reg[30] : (proc_35_data_FIFO_blk[30] | proc_35_data_PIPO_blk[30] | proc_35_start_FIFO_blk[30] | proc_35_TLF_FIFO_blk[30] | proc_35_input_sync_blk[30] | proc_35_output_sync_blk[30]);
    assign proc_35_data_FIFO_blk[31] = 1'b0;
    assign proc_35_data_PIPO_blk[31] = 1'b0;
    assign proc_35_start_FIFO_blk[31] = 1'b0;
    assign proc_35_TLF_FIFO_blk[31] = 1'b0;
    assign proc_35_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_35_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_35[31] = dl_detect_out ? proc_dep_vld_vec_35_reg[31] : (proc_35_data_FIFO_blk[31] | proc_35_data_PIPO_blk[31] | proc_35_start_FIFO_blk[31] | proc_35_TLF_FIFO_blk[31] | proc_35_input_sync_blk[31] | proc_35_output_sync_blk[31]);
    assign proc_35_data_FIFO_blk[32] = 1'b0;
    assign proc_35_data_PIPO_blk[32] = 1'b0;
    assign proc_35_start_FIFO_blk[32] = 1'b0;
    assign proc_35_TLF_FIFO_blk[32] = 1'b0;
    assign proc_35_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_30_U0_ap_ready & ProcessingElement_30_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_35_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_35[32] = dl_detect_out ? proc_dep_vld_vec_35_reg[32] : (proc_35_data_FIFO_blk[32] | proc_35_data_PIPO_blk[32] | proc_35_start_FIFO_blk[32] | proc_35_TLF_FIFO_blk[32] | proc_35_input_sync_blk[32] | proc_35_output_sync_blk[32]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_35_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_35_reg <= proc_dep_vld_vec_35;
        end
    end
    assign in_chan_dep_vld_vec_35[0] = dep_chan_vld_0_35;
    assign in_chan_dep_data_vec_35[39 : 0] = dep_chan_data_0_35;
    assign token_in_vec_35[0] = token_0_35;
    assign in_chan_dep_vld_vec_35[1] = dep_chan_vld_1_35;
    assign in_chan_dep_data_vec_35[79 : 40] = dep_chan_data_1_35;
    assign token_in_vec_35[1] = token_1_35;
    assign in_chan_dep_vld_vec_35[2] = dep_chan_vld_3_35;
    assign in_chan_dep_data_vec_35[119 : 80] = dep_chan_data_3_35;
    assign token_in_vec_35[2] = token_3_35;
    assign in_chan_dep_vld_vec_35[3] = dep_chan_vld_6_35;
    assign in_chan_dep_data_vec_35[159 : 120] = dep_chan_data_6_35;
    assign token_in_vec_35[3] = token_6_35;
    assign in_chan_dep_vld_vec_35[4] = dep_chan_vld_7_35;
    assign in_chan_dep_data_vec_35[199 : 160] = dep_chan_data_7_35;
    assign token_in_vec_35[4] = token_7_35;
    assign in_chan_dep_vld_vec_35[5] = dep_chan_vld_8_35;
    assign in_chan_dep_data_vec_35[239 : 200] = dep_chan_data_8_35;
    assign token_in_vec_35[5] = token_8_35;
    assign in_chan_dep_vld_vec_35[6] = dep_chan_vld_9_35;
    assign in_chan_dep_data_vec_35[279 : 240] = dep_chan_data_9_35;
    assign token_in_vec_35[6] = token_9_35;
    assign in_chan_dep_vld_vec_35[7] = dep_chan_vld_10_35;
    assign in_chan_dep_data_vec_35[319 : 280] = dep_chan_data_10_35;
    assign token_in_vec_35[7] = token_10_35;
    assign in_chan_dep_vld_vec_35[8] = dep_chan_vld_11_35;
    assign in_chan_dep_data_vec_35[359 : 320] = dep_chan_data_11_35;
    assign token_in_vec_35[8] = token_11_35;
    assign in_chan_dep_vld_vec_35[9] = dep_chan_vld_12_35;
    assign in_chan_dep_data_vec_35[399 : 360] = dep_chan_data_12_35;
    assign token_in_vec_35[9] = token_12_35;
    assign in_chan_dep_vld_vec_35[10] = dep_chan_vld_13_35;
    assign in_chan_dep_data_vec_35[439 : 400] = dep_chan_data_13_35;
    assign token_in_vec_35[10] = token_13_35;
    assign in_chan_dep_vld_vec_35[11] = dep_chan_vld_14_35;
    assign in_chan_dep_data_vec_35[479 : 440] = dep_chan_data_14_35;
    assign token_in_vec_35[11] = token_14_35;
    assign in_chan_dep_vld_vec_35[12] = dep_chan_vld_15_35;
    assign in_chan_dep_data_vec_35[519 : 480] = dep_chan_data_15_35;
    assign token_in_vec_35[12] = token_15_35;
    assign in_chan_dep_vld_vec_35[13] = dep_chan_vld_16_35;
    assign in_chan_dep_data_vec_35[559 : 520] = dep_chan_data_16_35;
    assign token_in_vec_35[13] = token_16_35;
    assign in_chan_dep_vld_vec_35[14] = dep_chan_vld_17_35;
    assign in_chan_dep_data_vec_35[599 : 560] = dep_chan_data_17_35;
    assign token_in_vec_35[14] = token_17_35;
    assign in_chan_dep_vld_vec_35[15] = dep_chan_vld_18_35;
    assign in_chan_dep_data_vec_35[639 : 600] = dep_chan_data_18_35;
    assign token_in_vec_35[15] = token_18_35;
    assign in_chan_dep_vld_vec_35[16] = dep_chan_vld_19_35;
    assign in_chan_dep_data_vec_35[679 : 640] = dep_chan_data_19_35;
    assign token_in_vec_35[16] = token_19_35;
    assign in_chan_dep_vld_vec_35[17] = dep_chan_vld_20_35;
    assign in_chan_dep_data_vec_35[719 : 680] = dep_chan_data_20_35;
    assign token_in_vec_35[17] = token_20_35;
    assign in_chan_dep_vld_vec_35[18] = dep_chan_vld_21_35;
    assign in_chan_dep_data_vec_35[759 : 720] = dep_chan_data_21_35;
    assign token_in_vec_35[18] = token_21_35;
    assign in_chan_dep_vld_vec_35[19] = dep_chan_vld_22_35;
    assign in_chan_dep_data_vec_35[799 : 760] = dep_chan_data_22_35;
    assign token_in_vec_35[19] = token_22_35;
    assign in_chan_dep_vld_vec_35[20] = dep_chan_vld_23_35;
    assign in_chan_dep_data_vec_35[839 : 800] = dep_chan_data_23_35;
    assign token_in_vec_35[20] = token_23_35;
    assign in_chan_dep_vld_vec_35[21] = dep_chan_vld_24_35;
    assign in_chan_dep_data_vec_35[879 : 840] = dep_chan_data_24_35;
    assign token_in_vec_35[21] = token_24_35;
    assign in_chan_dep_vld_vec_35[22] = dep_chan_vld_25_35;
    assign in_chan_dep_data_vec_35[919 : 880] = dep_chan_data_25_35;
    assign token_in_vec_35[22] = token_25_35;
    assign in_chan_dep_vld_vec_35[23] = dep_chan_vld_26_35;
    assign in_chan_dep_data_vec_35[959 : 920] = dep_chan_data_26_35;
    assign token_in_vec_35[23] = token_26_35;
    assign in_chan_dep_vld_vec_35[24] = dep_chan_vld_27_35;
    assign in_chan_dep_data_vec_35[999 : 960] = dep_chan_data_27_35;
    assign token_in_vec_35[24] = token_27_35;
    assign in_chan_dep_vld_vec_35[25] = dep_chan_vld_28_35;
    assign in_chan_dep_data_vec_35[1039 : 1000] = dep_chan_data_28_35;
    assign token_in_vec_35[25] = token_28_35;
    assign in_chan_dep_vld_vec_35[26] = dep_chan_vld_29_35;
    assign in_chan_dep_data_vec_35[1079 : 1040] = dep_chan_data_29_35;
    assign token_in_vec_35[26] = token_29_35;
    assign in_chan_dep_vld_vec_35[27] = dep_chan_vld_30_35;
    assign in_chan_dep_data_vec_35[1119 : 1080] = dep_chan_data_30_35;
    assign token_in_vec_35[27] = token_30_35;
    assign in_chan_dep_vld_vec_35[28] = dep_chan_vld_31_35;
    assign in_chan_dep_data_vec_35[1159 : 1120] = dep_chan_data_31_35;
    assign token_in_vec_35[28] = token_31_35;
    assign in_chan_dep_vld_vec_35[29] = dep_chan_vld_32_35;
    assign in_chan_dep_data_vec_35[1199 : 1160] = dep_chan_data_32_35;
    assign token_in_vec_35[29] = token_32_35;
    assign in_chan_dep_vld_vec_35[30] = dep_chan_vld_33_35;
    assign in_chan_dep_data_vec_35[1239 : 1200] = dep_chan_data_33_35;
    assign token_in_vec_35[30] = token_33_35;
    assign in_chan_dep_vld_vec_35[31] = dep_chan_vld_34_35;
    assign in_chan_dep_data_vec_35[1279 : 1240] = dep_chan_data_34_35;
    assign token_in_vec_35[31] = token_34_35;
    assign in_chan_dep_vld_vec_35[32] = dep_chan_vld_36_35;
    assign in_chan_dep_data_vec_35[1319 : 1280] = dep_chan_data_36_35;
    assign token_in_vec_35[32] = token_36_35;
    assign dep_chan_vld_35_34 = out_chan_dep_vld_vec_35[0];
    assign dep_chan_data_35_34 = out_chan_dep_data_35;
    assign token_35_34 = token_out_vec_35[0];
    assign dep_chan_vld_35_36 = out_chan_dep_vld_vec_35[1];
    assign dep_chan_data_35_36 = out_chan_dep_data_35;
    assign token_35_36 = token_out_vec_35[1];
    assign dep_chan_vld_35_0 = out_chan_dep_vld_vec_35[2];
    assign dep_chan_data_35_0 = out_chan_dep_data_35;
    assign token_35_0 = token_out_vec_35[2];
    assign dep_chan_vld_35_1 = out_chan_dep_vld_vec_35[3];
    assign dep_chan_data_35_1 = out_chan_dep_data_35;
    assign token_35_1 = token_out_vec_35[3];
    assign dep_chan_vld_35_3 = out_chan_dep_vld_vec_35[4];
    assign dep_chan_data_35_3 = out_chan_dep_data_35;
    assign token_35_3 = token_out_vec_35[4];
    assign dep_chan_vld_35_6 = out_chan_dep_vld_vec_35[5];
    assign dep_chan_data_35_6 = out_chan_dep_data_35;
    assign token_35_6 = token_out_vec_35[5];
    assign dep_chan_vld_35_7 = out_chan_dep_vld_vec_35[6];
    assign dep_chan_data_35_7 = out_chan_dep_data_35;
    assign token_35_7 = token_out_vec_35[6];
    assign dep_chan_vld_35_8 = out_chan_dep_vld_vec_35[7];
    assign dep_chan_data_35_8 = out_chan_dep_data_35;
    assign token_35_8 = token_out_vec_35[7];
    assign dep_chan_vld_35_9 = out_chan_dep_vld_vec_35[8];
    assign dep_chan_data_35_9 = out_chan_dep_data_35;
    assign token_35_9 = token_out_vec_35[8];
    assign dep_chan_vld_35_10 = out_chan_dep_vld_vec_35[9];
    assign dep_chan_data_35_10 = out_chan_dep_data_35;
    assign token_35_10 = token_out_vec_35[9];
    assign dep_chan_vld_35_11 = out_chan_dep_vld_vec_35[10];
    assign dep_chan_data_35_11 = out_chan_dep_data_35;
    assign token_35_11 = token_out_vec_35[10];
    assign dep_chan_vld_35_12 = out_chan_dep_vld_vec_35[11];
    assign dep_chan_data_35_12 = out_chan_dep_data_35;
    assign token_35_12 = token_out_vec_35[11];
    assign dep_chan_vld_35_13 = out_chan_dep_vld_vec_35[12];
    assign dep_chan_data_35_13 = out_chan_dep_data_35;
    assign token_35_13 = token_out_vec_35[12];
    assign dep_chan_vld_35_14 = out_chan_dep_vld_vec_35[13];
    assign dep_chan_data_35_14 = out_chan_dep_data_35;
    assign token_35_14 = token_out_vec_35[13];
    assign dep_chan_vld_35_15 = out_chan_dep_vld_vec_35[14];
    assign dep_chan_data_35_15 = out_chan_dep_data_35;
    assign token_35_15 = token_out_vec_35[14];
    assign dep_chan_vld_35_16 = out_chan_dep_vld_vec_35[15];
    assign dep_chan_data_35_16 = out_chan_dep_data_35;
    assign token_35_16 = token_out_vec_35[15];
    assign dep_chan_vld_35_17 = out_chan_dep_vld_vec_35[16];
    assign dep_chan_data_35_17 = out_chan_dep_data_35;
    assign token_35_17 = token_out_vec_35[16];
    assign dep_chan_vld_35_18 = out_chan_dep_vld_vec_35[17];
    assign dep_chan_data_35_18 = out_chan_dep_data_35;
    assign token_35_18 = token_out_vec_35[17];
    assign dep_chan_vld_35_19 = out_chan_dep_vld_vec_35[18];
    assign dep_chan_data_35_19 = out_chan_dep_data_35;
    assign token_35_19 = token_out_vec_35[18];
    assign dep_chan_vld_35_20 = out_chan_dep_vld_vec_35[19];
    assign dep_chan_data_35_20 = out_chan_dep_data_35;
    assign token_35_20 = token_out_vec_35[19];
    assign dep_chan_vld_35_21 = out_chan_dep_vld_vec_35[20];
    assign dep_chan_data_35_21 = out_chan_dep_data_35;
    assign token_35_21 = token_out_vec_35[20];
    assign dep_chan_vld_35_22 = out_chan_dep_vld_vec_35[21];
    assign dep_chan_data_35_22 = out_chan_dep_data_35;
    assign token_35_22 = token_out_vec_35[21];
    assign dep_chan_vld_35_23 = out_chan_dep_vld_vec_35[22];
    assign dep_chan_data_35_23 = out_chan_dep_data_35;
    assign token_35_23 = token_out_vec_35[22];
    assign dep_chan_vld_35_24 = out_chan_dep_vld_vec_35[23];
    assign dep_chan_data_35_24 = out_chan_dep_data_35;
    assign token_35_24 = token_out_vec_35[23];
    assign dep_chan_vld_35_25 = out_chan_dep_vld_vec_35[24];
    assign dep_chan_data_35_25 = out_chan_dep_data_35;
    assign token_35_25 = token_out_vec_35[24];
    assign dep_chan_vld_35_26 = out_chan_dep_vld_vec_35[25];
    assign dep_chan_data_35_26 = out_chan_dep_data_35;
    assign token_35_26 = token_out_vec_35[25];
    assign dep_chan_vld_35_27 = out_chan_dep_vld_vec_35[26];
    assign dep_chan_data_35_27 = out_chan_dep_data_35;
    assign token_35_27 = token_out_vec_35[26];
    assign dep_chan_vld_35_28 = out_chan_dep_vld_vec_35[27];
    assign dep_chan_data_35_28 = out_chan_dep_data_35;
    assign token_35_28 = token_out_vec_35[27];
    assign dep_chan_vld_35_29 = out_chan_dep_vld_vec_35[28];
    assign dep_chan_data_35_29 = out_chan_dep_data_35;
    assign token_35_29 = token_out_vec_35[28];
    assign dep_chan_vld_35_30 = out_chan_dep_vld_vec_35[29];
    assign dep_chan_data_35_30 = out_chan_dep_data_35;
    assign token_35_30 = token_out_vec_35[29];
    assign dep_chan_vld_35_31 = out_chan_dep_vld_vec_35[30];
    assign dep_chan_data_35_31 = out_chan_dep_data_35;
    assign token_35_31 = token_out_vec_35[30];
    assign dep_chan_vld_35_32 = out_chan_dep_vld_vec_35[31];
    assign dep_chan_data_35_32 = out_chan_dep_data_35;
    assign token_35_32 = token_out_vec_35[31];
    assign dep_chan_vld_35_33 = out_chan_dep_vld_vec_35[32];
    assign dep_chan_data_35_33 = out_chan_dep_data_35;
    assign token_35_33 = token_out_vec_35[32];

    // Process: ProcessingElement_31_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 36, 34, 34) MatrixMultiplicationKernel_hls_deadlock_detect_unit_36 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_36),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_36),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_36),
        .token_in_vec(token_in_vec_36),
        .dl_detect_in(dl_detect_out),
        .origin(origin[36]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_36),
        .out_chan_dep_data(out_chan_dep_data_36),
        .token_out_vec(token_out_vec_36),
        .dl_detect_out(dl_in_vec[36]));

    assign proc_36_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_190.aPipes_30_blk_n) | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_Pipeline_N_Pipeline_M_fu_199.bPipes_30_blk_n) | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_WriteC_Flattened_fu_221.cPipes_30_blk_n);
    assign proc_36_data_PIPO_blk[0] = 1'b0;
    assign proc_36_start_FIFO_blk[0] = 1'b0;
    assign proc_36_TLF_FIFO_blk[0] = 1'b0;
    assign proc_36_input_sync_blk[0] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_30_U0_ap_ready);
    assign proc_36_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_36[0] = dl_detect_out ? proc_dep_vld_vec_36_reg[0] : (proc_36_data_FIFO_blk[0] | proc_36_data_PIPO_blk[0] | proc_36_start_FIFO_blk[0] | proc_36_TLF_FIFO_blk[0] | proc_36_input_sync_blk[0] | proc_36_output_sync_blk[0]);
    assign proc_36_data_FIFO_blk[1] = 1'b0 | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_InitializeABuffer_Inner_InitializeABuffer_Outer_fu_190.aPipes_31_blk_n) | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_Pipeline_N_Pipeline_M_fu_199.bPipes_31_blk_n) | (~ProcessingElement_31_U0.grp_ProcessingElement_31_Pipeline_WriteC_Flattened_fu_221.cPipes_31_blk_n) | (~ProcessingElement_31_U0.size_n_c2_blk_n) | (~ProcessingElement_31_U0.size_k_c_blk_n) | (~ProcessingElement_31_U0.size_m_c10_blk_n);
    assign proc_36_data_PIPO_blk[1] = 1'b0;
    assign proc_36_start_FIFO_blk[1] = 1'b0 | (~start_for_ProcessingElement_U0_U.if_full_n & ProcessingElement_31_U0.ap_start & ~ProcessingElement_31_U0.real_start & (trans_in_cnt_3 == trans_out_cnt_3) & ~start_for_ProcessingElement_U0_U.if_read);
    assign proc_36_TLF_FIFO_blk[1] = 1'b0;
    assign proc_36_input_sync_blk[1] = 1'b0;
    assign proc_36_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_36[1] = dl_detect_out ? proc_dep_vld_vec_36_reg[1] : (proc_36_data_FIFO_blk[1] | proc_36_data_PIPO_blk[1] | proc_36_start_FIFO_blk[1] | proc_36_TLF_FIFO_blk[1] | proc_36_input_sync_blk[1] | proc_36_output_sync_blk[1]);
    assign proc_36_data_FIFO_blk[2] = 1'b0;
    assign proc_36_data_PIPO_blk[2] = 1'b0;
    assign proc_36_start_FIFO_blk[2] = 1'b0;
    assign proc_36_TLF_FIFO_blk[2] = 1'b0;
    assign proc_36_input_sync_blk[2] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_entry_proc_U0_ap_ready);
    assign proc_36_output_sync_blk[2] = 1'b0;
    assign proc_dep_vld_vec_36[2] = dl_detect_out ? proc_dep_vld_vec_36_reg[2] : (proc_36_data_FIFO_blk[2] | proc_36_data_PIPO_blk[2] | proc_36_start_FIFO_blk[2] | proc_36_TLF_FIFO_blk[2] | proc_36_input_sync_blk[2] | proc_36_output_sync_blk[2]);
    assign proc_36_data_FIFO_blk[3] = 1'b0;
    assign proc_36_data_PIPO_blk[3] = 1'b0;
    assign proc_36_start_FIFO_blk[3] = 1'b0;
    assign proc_36_TLF_FIFO_blk[3] = 1'b0;
    assign proc_36_input_sync_blk[3] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ReadA_U0_ap_ready);
    assign proc_36_output_sync_blk[3] = 1'b0;
    assign proc_dep_vld_vec_36[3] = dl_detect_out ? proc_dep_vld_vec_36_reg[3] : (proc_36_data_FIFO_blk[3] | proc_36_data_PIPO_blk[3] | proc_36_start_FIFO_blk[3] | proc_36_TLF_FIFO_blk[3] | proc_36_input_sync_blk[3] | proc_36_output_sync_blk[3]);
    assign proc_36_data_FIFO_blk[4] = 1'b0;
    assign proc_36_data_PIPO_blk[4] = 1'b0;
    assign proc_36_start_FIFO_blk[4] = 1'b0;
    assign proc_36_TLF_FIFO_blk[4] = 1'b0;
    assign proc_36_input_sync_blk[4] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ReadB_U0_ap_ready);
    assign proc_36_output_sync_blk[4] = 1'b0;
    assign proc_dep_vld_vec_36[4] = dl_detect_out ? proc_dep_vld_vec_36_reg[4] : (proc_36_data_FIFO_blk[4] | proc_36_data_PIPO_blk[4] | proc_36_start_FIFO_blk[4] | proc_36_TLF_FIFO_blk[4] | proc_36_input_sync_blk[4] | proc_36_output_sync_blk[4]);
    assign proc_36_data_FIFO_blk[5] = 1'b0;
    assign proc_36_data_PIPO_blk[5] = 1'b0;
    assign proc_36_start_FIFO_blk[5] = 1'b0;
    assign proc_36_TLF_FIFO_blk[5] = 1'b0;
    assign proc_36_input_sync_blk[5] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_1_U0_ap_ready);
    assign proc_36_output_sync_blk[5] = 1'b0;
    assign proc_dep_vld_vec_36[5] = dl_detect_out ? proc_dep_vld_vec_36_reg[5] : (proc_36_data_FIFO_blk[5] | proc_36_data_PIPO_blk[5] | proc_36_start_FIFO_blk[5] | proc_36_TLF_FIFO_blk[5] | proc_36_input_sync_blk[5] | proc_36_output_sync_blk[5]);
    assign proc_36_data_FIFO_blk[6] = 1'b0;
    assign proc_36_data_PIPO_blk[6] = 1'b0;
    assign proc_36_start_FIFO_blk[6] = 1'b0;
    assign proc_36_TLF_FIFO_blk[6] = 1'b0;
    assign proc_36_input_sync_blk[6] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_2_U0_ap_ready);
    assign proc_36_output_sync_blk[6] = 1'b0;
    assign proc_dep_vld_vec_36[6] = dl_detect_out ? proc_dep_vld_vec_36_reg[6] : (proc_36_data_FIFO_blk[6] | proc_36_data_PIPO_blk[6] | proc_36_start_FIFO_blk[6] | proc_36_TLF_FIFO_blk[6] | proc_36_input_sync_blk[6] | proc_36_output_sync_blk[6]);
    assign proc_36_data_FIFO_blk[7] = 1'b0;
    assign proc_36_data_PIPO_blk[7] = 1'b0;
    assign proc_36_start_FIFO_blk[7] = 1'b0;
    assign proc_36_TLF_FIFO_blk[7] = 1'b0;
    assign proc_36_input_sync_blk[7] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_3_U0_ap_ready);
    assign proc_36_output_sync_blk[7] = 1'b0;
    assign proc_dep_vld_vec_36[7] = dl_detect_out ? proc_dep_vld_vec_36_reg[7] : (proc_36_data_FIFO_blk[7] | proc_36_data_PIPO_blk[7] | proc_36_start_FIFO_blk[7] | proc_36_TLF_FIFO_blk[7] | proc_36_input_sync_blk[7] | proc_36_output_sync_blk[7]);
    assign proc_36_data_FIFO_blk[8] = 1'b0;
    assign proc_36_data_PIPO_blk[8] = 1'b0;
    assign proc_36_start_FIFO_blk[8] = 1'b0;
    assign proc_36_TLF_FIFO_blk[8] = 1'b0;
    assign proc_36_input_sync_blk[8] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_4_U0_ap_ready);
    assign proc_36_output_sync_blk[8] = 1'b0;
    assign proc_dep_vld_vec_36[8] = dl_detect_out ? proc_dep_vld_vec_36_reg[8] : (proc_36_data_FIFO_blk[8] | proc_36_data_PIPO_blk[8] | proc_36_start_FIFO_blk[8] | proc_36_TLF_FIFO_blk[8] | proc_36_input_sync_blk[8] | proc_36_output_sync_blk[8]);
    assign proc_36_data_FIFO_blk[9] = 1'b0;
    assign proc_36_data_PIPO_blk[9] = 1'b0;
    assign proc_36_start_FIFO_blk[9] = 1'b0;
    assign proc_36_TLF_FIFO_blk[9] = 1'b0;
    assign proc_36_input_sync_blk[9] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_5_U0_ap_ready);
    assign proc_36_output_sync_blk[9] = 1'b0;
    assign proc_dep_vld_vec_36[9] = dl_detect_out ? proc_dep_vld_vec_36_reg[9] : (proc_36_data_FIFO_blk[9] | proc_36_data_PIPO_blk[9] | proc_36_start_FIFO_blk[9] | proc_36_TLF_FIFO_blk[9] | proc_36_input_sync_blk[9] | proc_36_output_sync_blk[9]);
    assign proc_36_data_FIFO_blk[10] = 1'b0;
    assign proc_36_data_PIPO_blk[10] = 1'b0;
    assign proc_36_start_FIFO_blk[10] = 1'b0;
    assign proc_36_TLF_FIFO_blk[10] = 1'b0;
    assign proc_36_input_sync_blk[10] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_6_U0_ap_ready);
    assign proc_36_output_sync_blk[10] = 1'b0;
    assign proc_dep_vld_vec_36[10] = dl_detect_out ? proc_dep_vld_vec_36_reg[10] : (proc_36_data_FIFO_blk[10] | proc_36_data_PIPO_blk[10] | proc_36_start_FIFO_blk[10] | proc_36_TLF_FIFO_blk[10] | proc_36_input_sync_blk[10] | proc_36_output_sync_blk[10]);
    assign proc_36_data_FIFO_blk[11] = 1'b0;
    assign proc_36_data_PIPO_blk[11] = 1'b0;
    assign proc_36_start_FIFO_blk[11] = 1'b0;
    assign proc_36_TLF_FIFO_blk[11] = 1'b0;
    assign proc_36_input_sync_blk[11] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_7_U0_ap_ready);
    assign proc_36_output_sync_blk[11] = 1'b0;
    assign proc_dep_vld_vec_36[11] = dl_detect_out ? proc_dep_vld_vec_36_reg[11] : (proc_36_data_FIFO_blk[11] | proc_36_data_PIPO_blk[11] | proc_36_start_FIFO_blk[11] | proc_36_TLF_FIFO_blk[11] | proc_36_input_sync_blk[11] | proc_36_output_sync_blk[11]);
    assign proc_36_data_FIFO_blk[12] = 1'b0;
    assign proc_36_data_PIPO_blk[12] = 1'b0;
    assign proc_36_start_FIFO_blk[12] = 1'b0;
    assign proc_36_TLF_FIFO_blk[12] = 1'b0;
    assign proc_36_input_sync_blk[12] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_8_U0_ap_ready);
    assign proc_36_output_sync_blk[12] = 1'b0;
    assign proc_dep_vld_vec_36[12] = dl_detect_out ? proc_dep_vld_vec_36_reg[12] : (proc_36_data_FIFO_blk[12] | proc_36_data_PIPO_blk[12] | proc_36_start_FIFO_blk[12] | proc_36_TLF_FIFO_blk[12] | proc_36_input_sync_blk[12] | proc_36_output_sync_blk[12]);
    assign proc_36_data_FIFO_blk[13] = 1'b0;
    assign proc_36_data_PIPO_blk[13] = 1'b0;
    assign proc_36_start_FIFO_blk[13] = 1'b0;
    assign proc_36_TLF_FIFO_blk[13] = 1'b0;
    assign proc_36_input_sync_blk[13] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_9_U0_ap_ready);
    assign proc_36_output_sync_blk[13] = 1'b0;
    assign proc_dep_vld_vec_36[13] = dl_detect_out ? proc_dep_vld_vec_36_reg[13] : (proc_36_data_FIFO_blk[13] | proc_36_data_PIPO_blk[13] | proc_36_start_FIFO_blk[13] | proc_36_TLF_FIFO_blk[13] | proc_36_input_sync_blk[13] | proc_36_output_sync_blk[13]);
    assign proc_36_data_FIFO_blk[14] = 1'b0;
    assign proc_36_data_PIPO_blk[14] = 1'b0;
    assign proc_36_start_FIFO_blk[14] = 1'b0;
    assign proc_36_TLF_FIFO_blk[14] = 1'b0;
    assign proc_36_input_sync_blk[14] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_10_U0_ap_ready);
    assign proc_36_output_sync_blk[14] = 1'b0;
    assign proc_dep_vld_vec_36[14] = dl_detect_out ? proc_dep_vld_vec_36_reg[14] : (proc_36_data_FIFO_blk[14] | proc_36_data_PIPO_blk[14] | proc_36_start_FIFO_blk[14] | proc_36_TLF_FIFO_blk[14] | proc_36_input_sync_blk[14] | proc_36_output_sync_blk[14]);
    assign proc_36_data_FIFO_blk[15] = 1'b0;
    assign proc_36_data_PIPO_blk[15] = 1'b0;
    assign proc_36_start_FIFO_blk[15] = 1'b0;
    assign proc_36_TLF_FIFO_blk[15] = 1'b0;
    assign proc_36_input_sync_blk[15] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_11_U0_ap_ready);
    assign proc_36_output_sync_blk[15] = 1'b0;
    assign proc_dep_vld_vec_36[15] = dl_detect_out ? proc_dep_vld_vec_36_reg[15] : (proc_36_data_FIFO_blk[15] | proc_36_data_PIPO_blk[15] | proc_36_start_FIFO_blk[15] | proc_36_TLF_FIFO_blk[15] | proc_36_input_sync_blk[15] | proc_36_output_sync_blk[15]);
    assign proc_36_data_FIFO_blk[16] = 1'b0;
    assign proc_36_data_PIPO_blk[16] = 1'b0;
    assign proc_36_start_FIFO_blk[16] = 1'b0;
    assign proc_36_TLF_FIFO_blk[16] = 1'b0;
    assign proc_36_input_sync_blk[16] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_12_U0_ap_ready);
    assign proc_36_output_sync_blk[16] = 1'b0;
    assign proc_dep_vld_vec_36[16] = dl_detect_out ? proc_dep_vld_vec_36_reg[16] : (proc_36_data_FIFO_blk[16] | proc_36_data_PIPO_blk[16] | proc_36_start_FIFO_blk[16] | proc_36_TLF_FIFO_blk[16] | proc_36_input_sync_blk[16] | proc_36_output_sync_blk[16]);
    assign proc_36_data_FIFO_blk[17] = 1'b0;
    assign proc_36_data_PIPO_blk[17] = 1'b0;
    assign proc_36_start_FIFO_blk[17] = 1'b0;
    assign proc_36_TLF_FIFO_blk[17] = 1'b0;
    assign proc_36_input_sync_blk[17] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_13_U0_ap_ready);
    assign proc_36_output_sync_blk[17] = 1'b0;
    assign proc_dep_vld_vec_36[17] = dl_detect_out ? proc_dep_vld_vec_36_reg[17] : (proc_36_data_FIFO_blk[17] | proc_36_data_PIPO_blk[17] | proc_36_start_FIFO_blk[17] | proc_36_TLF_FIFO_blk[17] | proc_36_input_sync_blk[17] | proc_36_output_sync_blk[17]);
    assign proc_36_data_FIFO_blk[18] = 1'b0;
    assign proc_36_data_PIPO_blk[18] = 1'b0;
    assign proc_36_start_FIFO_blk[18] = 1'b0;
    assign proc_36_TLF_FIFO_blk[18] = 1'b0;
    assign proc_36_input_sync_blk[18] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_14_U0_ap_ready);
    assign proc_36_output_sync_blk[18] = 1'b0;
    assign proc_dep_vld_vec_36[18] = dl_detect_out ? proc_dep_vld_vec_36_reg[18] : (proc_36_data_FIFO_blk[18] | proc_36_data_PIPO_blk[18] | proc_36_start_FIFO_blk[18] | proc_36_TLF_FIFO_blk[18] | proc_36_input_sync_blk[18] | proc_36_output_sync_blk[18]);
    assign proc_36_data_FIFO_blk[19] = 1'b0;
    assign proc_36_data_PIPO_blk[19] = 1'b0;
    assign proc_36_start_FIFO_blk[19] = 1'b0;
    assign proc_36_TLF_FIFO_blk[19] = 1'b0;
    assign proc_36_input_sync_blk[19] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_15_U0_ap_ready);
    assign proc_36_output_sync_blk[19] = 1'b0;
    assign proc_dep_vld_vec_36[19] = dl_detect_out ? proc_dep_vld_vec_36_reg[19] : (proc_36_data_FIFO_blk[19] | proc_36_data_PIPO_blk[19] | proc_36_start_FIFO_blk[19] | proc_36_TLF_FIFO_blk[19] | proc_36_input_sync_blk[19] | proc_36_output_sync_blk[19]);
    assign proc_36_data_FIFO_blk[20] = 1'b0;
    assign proc_36_data_PIPO_blk[20] = 1'b0;
    assign proc_36_start_FIFO_blk[20] = 1'b0;
    assign proc_36_TLF_FIFO_blk[20] = 1'b0;
    assign proc_36_input_sync_blk[20] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_16_U0_ap_ready);
    assign proc_36_output_sync_blk[20] = 1'b0;
    assign proc_dep_vld_vec_36[20] = dl_detect_out ? proc_dep_vld_vec_36_reg[20] : (proc_36_data_FIFO_blk[20] | proc_36_data_PIPO_blk[20] | proc_36_start_FIFO_blk[20] | proc_36_TLF_FIFO_blk[20] | proc_36_input_sync_blk[20] | proc_36_output_sync_blk[20]);
    assign proc_36_data_FIFO_blk[21] = 1'b0;
    assign proc_36_data_PIPO_blk[21] = 1'b0;
    assign proc_36_start_FIFO_blk[21] = 1'b0;
    assign proc_36_TLF_FIFO_blk[21] = 1'b0;
    assign proc_36_input_sync_blk[21] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_17_U0_ap_ready);
    assign proc_36_output_sync_blk[21] = 1'b0;
    assign proc_dep_vld_vec_36[21] = dl_detect_out ? proc_dep_vld_vec_36_reg[21] : (proc_36_data_FIFO_blk[21] | proc_36_data_PIPO_blk[21] | proc_36_start_FIFO_blk[21] | proc_36_TLF_FIFO_blk[21] | proc_36_input_sync_blk[21] | proc_36_output_sync_blk[21]);
    assign proc_36_data_FIFO_blk[22] = 1'b0;
    assign proc_36_data_PIPO_blk[22] = 1'b0;
    assign proc_36_start_FIFO_blk[22] = 1'b0;
    assign proc_36_TLF_FIFO_blk[22] = 1'b0;
    assign proc_36_input_sync_blk[22] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_18_U0_ap_ready);
    assign proc_36_output_sync_blk[22] = 1'b0;
    assign proc_dep_vld_vec_36[22] = dl_detect_out ? proc_dep_vld_vec_36_reg[22] : (proc_36_data_FIFO_blk[22] | proc_36_data_PIPO_blk[22] | proc_36_start_FIFO_blk[22] | proc_36_TLF_FIFO_blk[22] | proc_36_input_sync_blk[22] | proc_36_output_sync_blk[22]);
    assign proc_36_data_FIFO_blk[23] = 1'b0;
    assign proc_36_data_PIPO_blk[23] = 1'b0;
    assign proc_36_start_FIFO_blk[23] = 1'b0;
    assign proc_36_TLF_FIFO_blk[23] = 1'b0;
    assign proc_36_input_sync_blk[23] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_19_U0_ap_ready);
    assign proc_36_output_sync_blk[23] = 1'b0;
    assign proc_dep_vld_vec_36[23] = dl_detect_out ? proc_dep_vld_vec_36_reg[23] : (proc_36_data_FIFO_blk[23] | proc_36_data_PIPO_blk[23] | proc_36_start_FIFO_blk[23] | proc_36_TLF_FIFO_blk[23] | proc_36_input_sync_blk[23] | proc_36_output_sync_blk[23]);
    assign proc_36_data_FIFO_blk[24] = 1'b0;
    assign proc_36_data_PIPO_blk[24] = 1'b0;
    assign proc_36_start_FIFO_blk[24] = 1'b0;
    assign proc_36_TLF_FIFO_blk[24] = 1'b0;
    assign proc_36_input_sync_blk[24] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_20_U0_ap_ready);
    assign proc_36_output_sync_blk[24] = 1'b0;
    assign proc_dep_vld_vec_36[24] = dl_detect_out ? proc_dep_vld_vec_36_reg[24] : (proc_36_data_FIFO_blk[24] | proc_36_data_PIPO_blk[24] | proc_36_start_FIFO_blk[24] | proc_36_TLF_FIFO_blk[24] | proc_36_input_sync_blk[24] | proc_36_output_sync_blk[24]);
    assign proc_36_data_FIFO_blk[25] = 1'b0;
    assign proc_36_data_PIPO_blk[25] = 1'b0;
    assign proc_36_start_FIFO_blk[25] = 1'b0;
    assign proc_36_TLF_FIFO_blk[25] = 1'b0;
    assign proc_36_input_sync_blk[25] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_21_U0_ap_ready);
    assign proc_36_output_sync_blk[25] = 1'b0;
    assign proc_dep_vld_vec_36[25] = dl_detect_out ? proc_dep_vld_vec_36_reg[25] : (proc_36_data_FIFO_blk[25] | proc_36_data_PIPO_blk[25] | proc_36_start_FIFO_blk[25] | proc_36_TLF_FIFO_blk[25] | proc_36_input_sync_blk[25] | proc_36_output_sync_blk[25]);
    assign proc_36_data_FIFO_blk[26] = 1'b0;
    assign proc_36_data_PIPO_blk[26] = 1'b0;
    assign proc_36_start_FIFO_blk[26] = 1'b0;
    assign proc_36_TLF_FIFO_blk[26] = 1'b0;
    assign proc_36_input_sync_blk[26] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_22_U0_ap_ready);
    assign proc_36_output_sync_blk[26] = 1'b0;
    assign proc_dep_vld_vec_36[26] = dl_detect_out ? proc_dep_vld_vec_36_reg[26] : (proc_36_data_FIFO_blk[26] | proc_36_data_PIPO_blk[26] | proc_36_start_FIFO_blk[26] | proc_36_TLF_FIFO_blk[26] | proc_36_input_sync_blk[26] | proc_36_output_sync_blk[26]);
    assign proc_36_data_FIFO_blk[27] = 1'b0;
    assign proc_36_data_PIPO_blk[27] = 1'b0;
    assign proc_36_start_FIFO_blk[27] = 1'b0;
    assign proc_36_TLF_FIFO_blk[27] = 1'b0;
    assign proc_36_input_sync_blk[27] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_23_U0_ap_ready);
    assign proc_36_output_sync_blk[27] = 1'b0;
    assign proc_dep_vld_vec_36[27] = dl_detect_out ? proc_dep_vld_vec_36_reg[27] : (proc_36_data_FIFO_blk[27] | proc_36_data_PIPO_blk[27] | proc_36_start_FIFO_blk[27] | proc_36_TLF_FIFO_blk[27] | proc_36_input_sync_blk[27] | proc_36_output_sync_blk[27]);
    assign proc_36_data_FIFO_blk[28] = 1'b0;
    assign proc_36_data_PIPO_blk[28] = 1'b0;
    assign proc_36_start_FIFO_blk[28] = 1'b0;
    assign proc_36_TLF_FIFO_blk[28] = 1'b0;
    assign proc_36_input_sync_blk[28] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_24_U0_ap_ready);
    assign proc_36_output_sync_blk[28] = 1'b0;
    assign proc_dep_vld_vec_36[28] = dl_detect_out ? proc_dep_vld_vec_36_reg[28] : (proc_36_data_FIFO_blk[28] | proc_36_data_PIPO_blk[28] | proc_36_start_FIFO_blk[28] | proc_36_TLF_FIFO_blk[28] | proc_36_input_sync_blk[28] | proc_36_output_sync_blk[28]);
    assign proc_36_data_FIFO_blk[29] = 1'b0;
    assign proc_36_data_PIPO_blk[29] = 1'b0;
    assign proc_36_start_FIFO_blk[29] = 1'b0;
    assign proc_36_TLF_FIFO_blk[29] = 1'b0;
    assign proc_36_input_sync_blk[29] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_25_U0_ap_ready);
    assign proc_36_output_sync_blk[29] = 1'b0;
    assign proc_dep_vld_vec_36[29] = dl_detect_out ? proc_dep_vld_vec_36_reg[29] : (proc_36_data_FIFO_blk[29] | proc_36_data_PIPO_blk[29] | proc_36_start_FIFO_blk[29] | proc_36_TLF_FIFO_blk[29] | proc_36_input_sync_blk[29] | proc_36_output_sync_blk[29]);
    assign proc_36_data_FIFO_blk[30] = 1'b0;
    assign proc_36_data_PIPO_blk[30] = 1'b0;
    assign proc_36_start_FIFO_blk[30] = 1'b0;
    assign proc_36_TLF_FIFO_blk[30] = 1'b0;
    assign proc_36_input_sync_blk[30] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_26_U0_ap_ready);
    assign proc_36_output_sync_blk[30] = 1'b0;
    assign proc_dep_vld_vec_36[30] = dl_detect_out ? proc_dep_vld_vec_36_reg[30] : (proc_36_data_FIFO_blk[30] | proc_36_data_PIPO_blk[30] | proc_36_start_FIFO_blk[30] | proc_36_TLF_FIFO_blk[30] | proc_36_input_sync_blk[30] | proc_36_output_sync_blk[30]);
    assign proc_36_data_FIFO_blk[31] = 1'b0;
    assign proc_36_data_PIPO_blk[31] = 1'b0;
    assign proc_36_start_FIFO_blk[31] = 1'b0;
    assign proc_36_TLF_FIFO_blk[31] = 1'b0;
    assign proc_36_input_sync_blk[31] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_27_U0_ap_ready);
    assign proc_36_output_sync_blk[31] = 1'b0;
    assign proc_dep_vld_vec_36[31] = dl_detect_out ? proc_dep_vld_vec_36_reg[31] : (proc_36_data_FIFO_blk[31] | proc_36_data_PIPO_blk[31] | proc_36_start_FIFO_blk[31] | proc_36_TLF_FIFO_blk[31] | proc_36_input_sync_blk[31] | proc_36_output_sync_blk[31]);
    assign proc_36_data_FIFO_blk[32] = 1'b0;
    assign proc_36_data_PIPO_blk[32] = 1'b0;
    assign proc_36_start_FIFO_blk[32] = 1'b0;
    assign proc_36_TLF_FIFO_blk[32] = 1'b0;
    assign proc_36_input_sync_blk[32] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_28_U0_ap_ready);
    assign proc_36_output_sync_blk[32] = 1'b0;
    assign proc_dep_vld_vec_36[32] = dl_detect_out ? proc_dep_vld_vec_36_reg[32] : (proc_36_data_FIFO_blk[32] | proc_36_data_PIPO_blk[32] | proc_36_start_FIFO_blk[32] | proc_36_TLF_FIFO_blk[32] | proc_36_input_sync_blk[32] | proc_36_output_sync_blk[32]);
    assign proc_36_data_FIFO_blk[33] = 1'b0;
    assign proc_36_data_PIPO_blk[33] = 1'b0;
    assign proc_36_start_FIFO_blk[33] = 1'b0;
    assign proc_36_TLF_FIFO_blk[33] = 1'b0;
    assign proc_36_input_sync_blk[33] = 1'b0 | (ap_sync_ProcessingElement_31_U0_ap_ready & ProcessingElement_31_U0.ap_idle & ~ap_sync_ProcessingElement_29_U0_ap_ready);
    assign proc_36_output_sync_blk[33] = 1'b0;
    assign proc_dep_vld_vec_36[33] = dl_detect_out ? proc_dep_vld_vec_36_reg[33] : (proc_36_data_FIFO_blk[33] | proc_36_data_PIPO_blk[33] | proc_36_start_FIFO_blk[33] | proc_36_TLF_FIFO_blk[33] | proc_36_input_sync_blk[33] | proc_36_output_sync_blk[33]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_36_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_36_reg <= proc_dep_vld_vec_36;
        end
    end
    assign in_chan_dep_vld_vec_36[0] = dep_chan_vld_0_36;
    assign in_chan_dep_data_vec_36[39 : 0] = dep_chan_data_0_36;
    assign token_in_vec_36[0] = token_0_36;
    assign in_chan_dep_vld_vec_36[1] = dep_chan_vld_1_36;
    assign in_chan_dep_data_vec_36[79 : 40] = dep_chan_data_1_36;
    assign token_in_vec_36[1] = token_1_36;
    assign in_chan_dep_vld_vec_36[2] = dep_chan_vld_3_36;
    assign in_chan_dep_data_vec_36[119 : 80] = dep_chan_data_3_36;
    assign token_in_vec_36[2] = token_3_36;
    assign in_chan_dep_vld_vec_36[3] = dep_chan_vld_6_36;
    assign in_chan_dep_data_vec_36[159 : 120] = dep_chan_data_6_36;
    assign token_in_vec_36[3] = token_6_36;
    assign in_chan_dep_vld_vec_36[4] = dep_chan_vld_7_36;
    assign in_chan_dep_data_vec_36[199 : 160] = dep_chan_data_7_36;
    assign token_in_vec_36[4] = token_7_36;
    assign in_chan_dep_vld_vec_36[5] = dep_chan_vld_8_36;
    assign in_chan_dep_data_vec_36[239 : 200] = dep_chan_data_8_36;
    assign token_in_vec_36[5] = token_8_36;
    assign in_chan_dep_vld_vec_36[6] = dep_chan_vld_9_36;
    assign in_chan_dep_data_vec_36[279 : 240] = dep_chan_data_9_36;
    assign token_in_vec_36[6] = token_9_36;
    assign in_chan_dep_vld_vec_36[7] = dep_chan_vld_10_36;
    assign in_chan_dep_data_vec_36[319 : 280] = dep_chan_data_10_36;
    assign token_in_vec_36[7] = token_10_36;
    assign in_chan_dep_vld_vec_36[8] = dep_chan_vld_11_36;
    assign in_chan_dep_data_vec_36[359 : 320] = dep_chan_data_11_36;
    assign token_in_vec_36[8] = token_11_36;
    assign in_chan_dep_vld_vec_36[9] = dep_chan_vld_12_36;
    assign in_chan_dep_data_vec_36[399 : 360] = dep_chan_data_12_36;
    assign token_in_vec_36[9] = token_12_36;
    assign in_chan_dep_vld_vec_36[10] = dep_chan_vld_13_36;
    assign in_chan_dep_data_vec_36[439 : 400] = dep_chan_data_13_36;
    assign token_in_vec_36[10] = token_13_36;
    assign in_chan_dep_vld_vec_36[11] = dep_chan_vld_14_36;
    assign in_chan_dep_data_vec_36[479 : 440] = dep_chan_data_14_36;
    assign token_in_vec_36[11] = token_14_36;
    assign in_chan_dep_vld_vec_36[12] = dep_chan_vld_15_36;
    assign in_chan_dep_data_vec_36[519 : 480] = dep_chan_data_15_36;
    assign token_in_vec_36[12] = token_15_36;
    assign in_chan_dep_vld_vec_36[13] = dep_chan_vld_16_36;
    assign in_chan_dep_data_vec_36[559 : 520] = dep_chan_data_16_36;
    assign token_in_vec_36[13] = token_16_36;
    assign in_chan_dep_vld_vec_36[14] = dep_chan_vld_17_36;
    assign in_chan_dep_data_vec_36[599 : 560] = dep_chan_data_17_36;
    assign token_in_vec_36[14] = token_17_36;
    assign in_chan_dep_vld_vec_36[15] = dep_chan_vld_18_36;
    assign in_chan_dep_data_vec_36[639 : 600] = dep_chan_data_18_36;
    assign token_in_vec_36[15] = token_18_36;
    assign in_chan_dep_vld_vec_36[16] = dep_chan_vld_19_36;
    assign in_chan_dep_data_vec_36[679 : 640] = dep_chan_data_19_36;
    assign token_in_vec_36[16] = token_19_36;
    assign in_chan_dep_vld_vec_36[17] = dep_chan_vld_20_36;
    assign in_chan_dep_data_vec_36[719 : 680] = dep_chan_data_20_36;
    assign token_in_vec_36[17] = token_20_36;
    assign in_chan_dep_vld_vec_36[18] = dep_chan_vld_21_36;
    assign in_chan_dep_data_vec_36[759 : 720] = dep_chan_data_21_36;
    assign token_in_vec_36[18] = token_21_36;
    assign in_chan_dep_vld_vec_36[19] = dep_chan_vld_22_36;
    assign in_chan_dep_data_vec_36[799 : 760] = dep_chan_data_22_36;
    assign token_in_vec_36[19] = token_22_36;
    assign in_chan_dep_vld_vec_36[20] = dep_chan_vld_23_36;
    assign in_chan_dep_data_vec_36[839 : 800] = dep_chan_data_23_36;
    assign token_in_vec_36[20] = token_23_36;
    assign in_chan_dep_vld_vec_36[21] = dep_chan_vld_24_36;
    assign in_chan_dep_data_vec_36[879 : 840] = dep_chan_data_24_36;
    assign token_in_vec_36[21] = token_24_36;
    assign in_chan_dep_vld_vec_36[22] = dep_chan_vld_25_36;
    assign in_chan_dep_data_vec_36[919 : 880] = dep_chan_data_25_36;
    assign token_in_vec_36[22] = token_25_36;
    assign in_chan_dep_vld_vec_36[23] = dep_chan_vld_26_36;
    assign in_chan_dep_data_vec_36[959 : 920] = dep_chan_data_26_36;
    assign token_in_vec_36[23] = token_26_36;
    assign in_chan_dep_vld_vec_36[24] = dep_chan_vld_27_36;
    assign in_chan_dep_data_vec_36[999 : 960] = dep_chan_data_27_36;
    assign token_in_vec_36[24] = token_27_36;
    assign in_chan_dep_vld_vec_36[25] = dep_chan_vld_28_36;
    assign in_chan_dep_data_vec_36[1039 : 1000] = dep_chan_data_28_36;
    assign token_in_vec_36[25] = token_28_36;
    assign in_chan_dep_vld_vec_36[26] = dep_chan_vld_29_36;
    assign in_chan_dep_data_vec_36[1079 : 1040] = dep_chan_data_29_36;
    assign token_in_vec_36[26] = token_29_36;
    assign in_chan_dep_vld_vec_36[27] = dep_chan_vld_30_36;
    assign in_chan_dep_data_vec_36[1119 : 1080] = dep_chan_data_30_36;
    assign token_in_vec_36[27] = token_30_36;
    assign in_chan_dep_vld_vec_36[28] = dep_chan_vld_31_36;
    assign in_chan_dep_data_vec_36[1159 : 1120] = dep_chan_data_31_36;
    assign token_in_vec_36[28] = token_31_36;
    assign in_chan_dep_vld_vec_36[29] = dep_chan_vld_32_36;
    assign in_chan_dep_data_vec_36[1199 : 1160] = dep_chan_data_32_36;
    assign token_in_vec_36[29] = token_32_36;
    assign in_chan_dep_vld_vec_36[30] = dep_chan_vld_33_36;
    assign in_chan_dep_data_vec_36[1239 : 1200] = dep_chan_data_33_36;
    assign token_in_vec_36[30] = token_33_36;
    assign in_chan_dep_vld_vec_36[31] = dep_chan_vld_34_36;
    assign in_chan_dep_data_vec_36[1279 : 1240] = dep_chan_data_34_36;
    assign token_in_vec_36[31] = token_34_36;
    assign in_chan_dep_vld_vec_36[32] = dep_chan_vld_35_36;
    assign in_chan_dep_data_vec_36[1319 : 1280] = dep_chan_data_35_36;
    assign token_in_vec_36[32] = token_35_36;
    assign in_chan_dep_vld_vec_36[33] = dep_chan_vld_37_36;
    assign in_chan_dep_data_vec_36[1359 : 1320] = dep_chan_data_37_36;
    assign token_in_vec_36[33] = token_37_36;
    assign dep_chan_vld_36_35 = out_chan_dep_vld_vec_36[0];
    assign dep_chan_data_36_35 = out_chan_dep_data_36;
    assign token_36_35 = token_out_vec_36[0];
    assign dep_chan_vld_36_37 = out_chan_dep_vld_vec_36[1];
    assign dep_chan_data_36_37 = out_chan_dep_data_36;
    assign token_36_37 = token_out_vec_36[1];
    assign dep_chan_vld_36_0 = out_chan_dep_vld_vec_36[2];
    assign dep_chan_data_36_0 = out_chan_dep_data_36;
    assign token_36_0 = token_out_vec_36[2];
    assign dep_chan_vld_36_1 = out_chan_dep_vld_vec_36[3];
    assign dep_chan_data_36_1 = out_chan_dep_data_36;
    assign token_36_1 = token_out_vec_36[3];
    assign dep_chan_vld_36_3 = out_chan_dep_vld_vec_36[4];
    assign dep_chan_data_36_3 = out_chan_dep_data_36;
    assign token_36_3 = token_out_vec_36[4];
    assign dep_chan_vld_36_6 = out_chan_dep_vld_vec_36[5];
    assign dep_chan_data_36_6 = out_chan_dep_data_36;
    assign token_36_6 = token_out_vec_36[5];
    assign dep_chan_vld_36_7 = out_chan_dep_vld_vec_36[6];
    assign dep_chan_data_36_7 = out_chan_dep_data_36;
    assign token_36_7 = token_out_vec_36[6];
    assign dep_chan_vld_36_8 = out_chan_dep_vld_vec_36[7];
    assign dep_chan_data_36_8 = out_chan_dep_data_36;
    assign token_36_8 = token_out_vec_36[7];
    assign dep_chan_vld_36_9 = out_chan_dep_vld_vec_36[8];
    assign dep_chan_data_36_9 = out_chan_dep_data_36;
    assign token_36_9 = token_out_vec_36[8];
    assign dep_chan_vld_36_10 = out_chan_dep_vld_vec_36[9];
    assign dep_chan_data_36_10 = out_chan_dep_data_36;
    assign token_36_10 = token_out_vec_36[9];
    assign dep_chan_vld_36_11 = out_chan_dep_vld_vec_36[10];
    assign dep_chan_data_36_11 = out_chan_dep_data_36;
    assign token_36_11 = token_out_vec_36[10];
    assign dep_chan_vld_36_12 = out_chan_dep_vld_vec_36[11];
    assign dep_chan_data_36_12 = out_chan_dep_data_36;
    assign token_36_12 = token_out_vec_36[11];
    assign dep_chan_vld_36_13 = out_chan_dep_vld_vec_36[12];
    assign dep_chan_data_36_13 = out_chan_dep_data_36;
    assign token_36_13 = token_out_vec_36[12];
    assign dep_chan_vld_36_14 = out_chan_dep_vld_vec_36[13];
    assign dep_chan_data_36_14 = out_chan_dep_data_36;
    assign token_36_14 = token_out_vec_36[13];
    assign dep_chan_vld_36_15 = out_chan_dep_vld_vec_36[14];
    assign dep_chan_data_36_15 = out_chan_dep_data_36;
    assign token_36_15 = token_out_vec_36[14];
    assign dep_chan_vld_36_16 = out_chan_dep_vld_vec_36[15];
    assign dep_chan_data_36_16 = out_chan_dep_data_36;
    assign token_36_16 = token_out_vec_36[15];
    assign dep_chan_vld_36_17 = out_chan_dep_vld_vec_36[16];
    assign dep_chan_data_36_17 = out_chan_dep_data_36;
    assign token_36_17 = token_out_vec_36[16];
    assign dep_chan_vld_36_18 = out_chan_dep_vld_vec_36[17];
    assign dep_chan_data_36_18 = out_chan_dep_data_36;
    assign token_36_18 = token_out_vec_36[17];
    assign dep_chan_vld_36_19 = out_chan_dep_vld_vec_36[18];
    assign dep_chan_data_36_19 = out_chan_dep_data_36;
    assign token_36_19 = token_out_vec_36[18];
    assign dep_chan_vld_36_20 = out_chan_dep_vld_vec_36[19];
    assign dep_chan_data_36_20 = out_chan_dep_data_36;
    assign token_36_20 = token_out_vec_36[19];
    assign dep_chan_vld_36_21 = out_chan_dep_vld_vec_36[20];
    assign dep_chan_data_36_21 = out_chan_dep_data_36;
    assign token_36_21 = token_out_vec_36[20];
    assign dep_chan_vld_36_22 = out_chan_dep_vld_vec_36[21];
    assign dep_chan_data_36_22 = out_chan_dep_data_36;
    assign token_36_22 = token_out_vec_36[21];
    assign dep_chan_vld_36_23 = out_chan_dep_vld_vec_36[22];
    assign dep_chan_data_36_23 = out_chan_dep_data_36;
    assign token_36_23 = token_out_vec_36[22];
    assign dep_chan_vld_36_24 = out_chan_dep_vld_vec_36[23];
    assign dep_chan_data_36_24 = out_chan_dep_data_36;
    assign token_36_24 = token_out_vec_36[23];
    assign dep_chan_vld_36_25 = out_chan_dep_vld_vec_36[24];
    assign dep_chan_data_36_25 = out_chan_dep_data_36;
    assign token_36_25 = token_out_vec_36[24];
    assign dep_chan_vld_36_26 = out_chan_dep_vld_vec_36[25];
    assign dep_chan_data_36_26 = out_chan_dep_data_36;
    assign token_36_26 = token_out_vec_36[25];
    assign dep_chan_vld_36_27 = out_chan_dep_vld_vec_36[26];
    assign dep_chan_data_36_27 = out_chan_dep_data_36;
    assign token_36_27 = token_out_vec_36[26];
    assign dep_chan_vld_36_28 = out_chan_dep_vld_vec_36[27];
    assign dep_chan_data_36_28 = out_chan_dep_data_36;
    assign token_36_28 = token_out_vec_36[27];
    assign dep_chan_vld_36_29 = out_chan_dep_vld_vec_36[28];
    assign dep_chan_data_36_29 = out_chan_dep_data_36;
    assign token_36_29 = token_out_vec_36[28];
    assign dep_chan_vld_36_30 = out_chan_dep_vld_vec_36[29];
    assign dep_chan_data_36_30 = out_chan_dep_data_36;
    assign token_36_30 = token_out_vec_36[29];
    assign dep_chan_vld_36_31 = out_chan_dep_vld_vec_36[30];
    assign dep_chan_data_36_31 = out_chan_dep_data_36;
    assign token_36_31 = token_out_vec_36[30];
    assign dep_chan_vld_36_32 = out_chan_dep_vld_vec_36[31];
    assign dep_chan_data_36_32 = out_chan_dep_data_36;
    assign token_36_32 = token_out_vec_36[31];
    assign dep_chan_vld_36_33 = out_chan_dep_vld_vec_36[32];
    assign dep_chan_data_36_33 = out_chan_dep_data_36;
    assign token_36_33 = token_out_vec_36[32];
    assign dep_chan_vld_36_34 = out_chan_dep_vld_vec_36[33];
    assign dep_chan_data_36_34 = out_chan_dep_data_36;
    assign token_36_34 = token_out_vec_36[33];

    // Process: ProcessingElement_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 37, 2, 2) MatrixMultiplicationKernel_hls_deadlock_detect_unit_37 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_37),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_37),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_37),
        .token_in_vec(token_in_vec_37),
        .dl_detect_in(dl_detect_out),
        .origin(origin[37]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_37),
        .out_chan_dep_data(out_chan_dep_data_37),
        .token_out_vec(token_out_vec_37),
        .dl_detect_out(dl_in_vec[37]));

    assign proc_37_data_FIFO_blk[0] = 1'b0 | (~ProcessingElement_U0.grp_ProcessingElement_Pipeline_Pipeline_N_Pipeline_M_fu_159.aPipes_31_blk_n) | (~ProcessingElement_U0.grp_ProcessingElement_Pipeline_Pipeline_N_Pipeline_M_fu_159.bPipes_31_blk_n) | (~ProcessingElement_U0.grp_ProcessingElement_Pipeline_WriteC_Flattened_fu_177.cPipes_31_blk_n) | (~ProcessingElement_U0.size_n_blk_n) | (~ProcessingElement_U0.size_k_blk_n) | (~ProcessingElement_U0.size_m_blk_n);
    assign proc_37_data_PIPO_blk[0] = 1'b0;
    assign proc_37_start_FIFO_blk[0] = 1'b0 | (~start_for_ProcessingElement_U0_U.if_empty_n & ProcessingElement_U0.ap_idle & ~start_for_ProcessingElement_U0_U.if_write);
    assign proc_37_TLF_FIFO_blk[0] = 1'b0;
    assign proc_37_input_sync_blk[0] = 1'b0;
    assign proc_37_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_37[0] = dl_detect_out ? proc_dep_vld_vec_37_reg[0] : (proc_37_data_FIFO_blk[0] | proc_37_data_PIPO_blk[0] | proc_37_start_FIFO_blk[0] | proc_37_TLF_FIFO_blk[0] | proc_37_input_sync_blk[0] | proc_37_output_sync_blk[0]);
    assign proc_37_data_FIFO_blk[1] = 1'b0;
    assign proc_37_data_PIPO_blk[1] = 1'b0;
    assign proc_37_start_FIFO_blk[1] = 1'b0;
    assign proc_37_TLF_FIFO_blk[1] = 1'b0;
    assign proc_37_input_sync_blk[1] = 1'b0;
    assign proc_37_output_sync_blk[1] = 1'b0 | (ap_done_reg_0 & ProcessingElement_U0.ap_done & ~WriteC_U0.ap_done);
    assign proc_dep_vld_vec_37[1] = dl_detect_out ? proc_dep_vld_vec_37_reg[1] : (proc_37_data_FIFO_blk[1] | proc_37_data_PIPO_blk[1] | proc_37_start_FIFO_blk[1] | proc_37_TLF_FIFO_blk[1] | proc_37_input_sync_blk[1] | proc_37_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_37_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_37_reg <= proc_dep_vld_vec_37;
        end
    end
    assign in_chan_dep_vld_vec_37[0] = dep_chan_vld_36_37;
    assign in_chan_dep_data_vec_37[39 : 0] = dep_chan_data_36_37;
    assign token_in_vec_37[0] = token_36_37;
    assign in_chan_dep_vld_vec_37[1] = dep_chan_vld_39_37;
    assign in_chan_dep_data_vec_37[79 : 40] = dep_chan_data_39_37;
    assign token_in_vec_37[1] = token_39_37;
    assign dep_chan_vld_37_36 = out_chan_dep_vld_vec_37[0];
    assign dep_chan_data_37_36 = out_chan_dep_data_37;
    assign token_37_36 = token_out_vec_37[0];
    assign dep_chan_vld_37_39 = out_chan_dep_vld_vec_37[1];
    assign dep_chan_data_37_39 = out_chan_dep_data_37;
    assign token_37_39 = token_out_vec_37[1];

    // Process: ConvertWidthC_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 38, 2, 2) MatrixMultiplicationKernel_hls_deadlock_detect_unit_38 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_38),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_38),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_38),
        .token_in_vec(token_in_vec_38),
        .dl_detect_in(dl_detect_out),
        .origin(origin[38]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_38),
        .out_chan_dep_data(out_chan_dep_data_38),
        .token_out_vec(token_out_vec_38),
        .dl_detect_out(dl_in_vec[38]));

    assign proc_38_data_FIFO_blk[0] = 1'b0 | (~ConvertWidthC_U0.grp_ConvertWidthC_Pipeline_ConvertWidthC_N_ConvertWidthC_M_VITIS_LOOP_339_1_fu_84.cPipes_0_blk_n) | (~ConvertWidthC_U0.size_n_blk_n) | (~ConvertWidthC_U0.size_m_blk_n);
    assign proc_38_data_PIPO_blk[0] = 1'b0;
    assign proc_38_start_FIFO_blk[0] = 1'b0 | (~start_for_ConvertWidthC_U0_U.if_empty_n & ConvertWidthC_U0.ap_idle & ~start_for_ConvertWidthC_U0_U.if_write);
    assign proc_38_TLF_FIFO_blk[0] = 1'b0;
    assign proc_38_input_sync_blk[0] = 1'b0;
    assign proc_38_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_38[0] = dl_detect_out ? proc_dep_vld_vec_38_reg[0] : (proc_38_data_FIFO_blk[0] | proc_38_data_PIPO_blk[0] | proc_38_start_FIFO_blk[0] | proc_38_TLF_FIFO_blk[0] | proc_38_input_sync_blk[0] | proc_38_output_sync_blk[0]);
    assign proc_38_data_FIFO_blk[1] = 1'b0 | (~ConvertWidthC_U0.grp_ConvertWidthC_Pipeline_ConvertWidthC_N_ConvertWidthC_M_VITIS_LOOP_339_1_fu_84.cMemory_blk_n) | (~ConvertWidthC_U0.size_n_c_blk_n) | (~ConvertWidthC_U0.size_m_c_blk_n);
    assign proc_38_data_PIPO_blk[1] = 1'b0;
    assign proc_38_start_FIFO_blk[1] = 1'b0;
    assign proc_38_TLF_FIFO_blk[1] = 1'b0;
    assign proc_38_input_sync_blk[1] = 1'b0;
    assign proc_38_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_38[1] = dl_detect_out ? proc_dep_vld_vec_38_reg[1] : (proc_38_data_FIFO_blk[1] | proc_38_data_PIPO_blk[1] | proc_38_start_FIFO_blk[1] | proc_38_TLF_FIFO_blk[1] | proc_38_input_sync_blk[1] | proc_38_output_sync_blk[1]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_38_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_38_reg <= proc_dep_vld_vec_38;
        end
    end
    assign in_chan_dep_vld_vec_38[0] = dep_chan_vld_6_38;
    assign in_chan_dep_data_vec_38[39 : 0] = dep_chan_data_6_38;
    assign token_in_vec_38[0] = token_6_38;
    assign in_chan_dep_vld_vec_38[1] = dep_chan_vld_39_38;
    assign in_chan_dep_data_vec_38[79 : 40] = dep_chan_data_39_38;
    assign token_in_vec_38[1] = token_39_38;
    assign dep_chan_vld_38_6 = out_chan_dep_vld_vec_38[0];
    assign dep_chan_data_38_6 = out_chan_dep_data_38;
    assign token_38_6 = token_out_vec_38[0];
    assign dep_chan_vld_38_39 = out_chan_dep_vld_vec_38[1];
    assign dep_chan_data_38_39 = out_chan_dep_data_38;
    assign token_38_39 = token_out_vec_38[1];

    // Process: WriteC_U0
    MatrixMultiplicationKernel_hls_deadlock_detect_unit #(40, 39, 3, 3) MatrixMultiplicationKernel_hls_deadlock_detect_unit_39 (
        .reset(dl_reset),
        .clock(dl_clock),
        .proc_dep_vld_vec(proc_dep_vld_vec_39),
        .in_chan_dep_vld_vec(in_chan_dep_vld_vec_39),
        .in_chan_dep_data_vec(in_chan_dep_data_vec_39),
        .token_in_vec(token_in_vec_39),
        .dl_detect_in(dl_detect_out),
        .origin(origin[39]),
        .token_clear(token_clear),
        .out_chan_dep_vld_vec(out_chan_dep_vld_vec_39),
        .out_chan_dep_data(out_chan_dep_data_39),
        .token_out_vec(token_out_vec_39),
        .dl_detect_out(dl_in_vec[39]));

    assign proc_39_data_FIFO_blk[0] = 1'b0 | (~WriteC_U0.grp_WriteC_Pipeline_WriteC_OuterTile_N_WriteC_OuterTile_M_WriteC_N1_WriteC_M1_fu_82.cMemory_blk_n) | (~WriteC_U0.size_n_blk_n) | (~WriteC_U0.size_m_blk_n);
    assign proc_39_data_PIPO_blk[0] = 1'b0;
    assign proc_39_start_FIFO_blk[0] = 1'b0;
    assign proc_39_TLF_FIFO_blk[0] = 1'b0;
    assign proc_39_input_sync_blk[0] = 1'b0;
    assign proc_39_output_sync_blk[0] = 1'b0;
    assign proc_dep_vld_vec_39[0] = dl_detect_out ? proc_dep_vld_vec_39_reg[0] : (proc_39_data_FIFO_blk[0] | proc_39_data_PIPO_blk[0] | proc_39_start_FIFO_blk[0] | proc_39_TLF_FIFO_blk[0] | proc_39_input_sync_blk[0] | proc_39_output_sync_blk[0]);
    assign proc_39_data_FIFO_blk[1] = 1'b0 | (~WriteC_U0.memory_blk_n);
    assign proc_39_data_PIPO_blk[1] = 1'b0;
    assign proc_39_start_FIFO_blk[1] = 1'b0 | (~start_for_WriteC_U0_U.if_empty_n & WriteC_U0.ap_idle & ~start_for_WriteC_U0_U.if_write);
    assign proc_39_TLF_FIFO_blk[1] = 1'b0;
    assign proc_39_input_sync_blk[1] = 1'b0;
    assign proc_39_output_sync_blk[1] = 1'b0;
    assign proc_dep_vld_vec_39[1] = dl_detect_out ? proc_dep_vld_vec_39_reg[1] : (proc_39_data_FIFO_blk[1] | proc_39_data_PIPO_blk[1] | proc_39_start_FIFO_blk[1] | proc_39_TLF_FIFO_blk[1] | proc_39_input_sync_blk[1] | proc_39_output_sync_blk[1]);
    assign proc_39_data_FIFO_blk[2] = 1'b0;
    assign proc_39_data_PIPO_blk[2] = 1'b0;
    assign proc_39_start_FIFO_blk[2] = 1'b0;
    assign proc_39_TLF_FIFO_blk[2] = 1'b0;
    assign proc_39_input_sync_blk[2] = 1'b0;
    assign proc_39_output_sync_blk[2] = 1'b0 | (ap_done_reg_1 & WriteC_U0.ap_done & ~ProcessingElement_U0.ap_done);
    assign proc_dep_vld_vec_39[2] = dl_detect_out ? proc_dep_vld_vec_39_reg[2] : (proc_39_data_FIFO_blk[2] | proc_39_data_PIPO_blk[2] | proc_39_start_FIFO_blk[2] | proc_39_TLF_FIFO_blk[2] | proc_39_input_sync_blk[2] | proc_39_output_sync_blk[2]);
    always @ (negedge dl_reset or posedge dl_clock) begin
        if (~dl_reset) begin
            proc_dep_vld_vec_39_reg <= 'b0;
        end
        else begin
            proc_dep_vld_vec_39_reg <= proc_dep_vld_vec_39;
        end
    end
    assign in_chan_dep_vld_vec_39[0] = dep_chan_vld_0_39;
    assign in_chan_dep_data_vec_39[39 : 0] = dep_chan_data_0_39;
    assign token_in_vec_39[0] = token_0_39;
    assign in_chan_dep_vld_vec_39[1] = dep_chan_vld_37_39;
    assign in_chan_dep_data_vec_39[79 : 40] = dep_chan_data_37_39;
    assign token_in_vec_39[1] = token_37_39;
    assign in_chan_dep_vld_vec_39[2] = dep_chan_vld_38_39;
    assign in_chan_dep_data_vec_39[119 : 80] = dep_chan_data_38_39;
    assign token_in_vec_39[2] = token_38_39;
    assign dep_chan_vld_39_38 = out_chan_dep_vld_vec_39[0];
    assign dep_chan_data_39_38 = out_chan_dep_data_39;
    assign token_39_38 = token_out_vec_39[0];
    assign dep_chan_vld_39_0 = out_chan_dep_vld_vec_39[1];
    assign dep_chan_data_39_0 = out_chan_dep_data_39;
    assign token_39_0 = token_out_vec_39[1];
    assign dep_chan_vld_39_37 = out_chan_dep_vld_vec_39[2];
    assign dep_chan_data_39_37 = out_chan_dep_data_39;
    assign token_39_37 = token_out_vec_39[2];


`include "MatrixMultiplicationKernel_hls_deadlock_report_unit.vh"
